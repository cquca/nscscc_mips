`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hmgGeiuU85OrkJlied/6OZ/LeCurFTEBnHiOPfVoXA+EBs+SHGB41VJIX4wobZy/n6y6FSxdzhAI
UKc9ut4Wnw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
S32LRXMx8RCmugnJlaKzfXlJUfIoaCF0uAe00huNbMYEr70MUEkXTAEuGHUdTsq+Y7V7DDN+ruip
JFkAzXZl//RBL4IS2hjGrLOBq7LOXcEgWjZMikYvYnGMBRDHX1ezkLjxJz1F5v9yzKInXQAxdpND
jzmSV87ClNMFvpUYjR8=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Oe47XaGVPilIcDcNRpYdlMIAuesZfXMx5o6OCMqxqSsHA7G7my7ZlpgyH6sg+WO4mMr2hv5ufFSE
ybEmiT0drndcQq14JQFKsuqEBBByNiNzyZMHin3AvnOfcXuC+acQUJ7nkEM8HBFdEBujyh7peq5T
WCYfwZknQvvgrbPdCVE=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AejPo+ecBHd1+UuTZ9CZcLDWKbgTnq/yjgV3bZNYSdJN9ZqjS5dNOpCZjMZkaKeSNurvkmv3btwN
QCoQ8KQvstc9H1xBUobbP3XTMj/v3SbShQUihj5HyhrtGcv5zK2fSTSNosOZXnvAqr5VpFw+aBPQ
E9glw4zbZUN6pb67AhW+2ojsvG4JUBg7+czW9pu2F/WJ1FSi6yVeQV1TjNWm3W9q35f4t4ypylmd
6t+6F/6w6p45f76ABuvu1L4ATGL1IwteKDYqTbCIZ2mdfK5/JpEqLUOUtTkPBqERB47tGCzL1BNl
aWPn0U4VZ7wFvMlREA+2i1d31m7bt16jzHyXqg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
etNUku/cmg58IjND4HdAEtq4g9P5gsK2GDk0V2TyNr6r4RUBxzZtzO5wWJ3k0nFu0iMR/taAl/q3
XxSMhdwgMRXHLr3FoWHRvuzGFsFUu96TB7+5yQl7g6kG1xbdq1J2Q69tS2BY52VjSagkxOGqOrIs
xs9rF7lQbqoFJmPDw23FADAiEy1/8YQ0P9vtk9kYt82E6YqR+CLUGCaYRf+GdyAaRpaacsy/voG6
xxPfQC0TMMZQl7pBvtex8slqAQJduzwXQoPdGykBon+GEX567ajGEK4eF+G3fWKaAeMEppi8AF/3
MwdCPcWFYo1/nrHqqtuq+BfbpEQdSHreQTDEJg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Qwac+t8oNxRmBVPNv19fdihUJ5FSXsBxRWk6ZZT6YpVoz5Hz9p3SclbEBb5hxqg+5rd0yG0zlJ4s
oe5zk3qs9ka4O6UWoAT4v1Avo9dyxVqOLgKd4uZ7tuuILBJE+H+GJ3puSWInbDNeX+xhkSUfd0Ou
dSgPEtW59ZYGfvxVhjLwMS813lJTrx6GPwFPmAwomNuV6eZEB1DDWA1F7ea5yYKw9hMT6SVyC7tF
g+dJfum0hU5Dsw1myNuVtay8j/OOfTRgZ8nkXe9HKwrvXfWHy39J1FGpTDKlztl2AcS+iRh2nk/S
04zDeLNWUrVHGb8SZgjBE99o2MEsWa0O0okSUA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11005744)
`protect data_block
b8i9C4PHAWDHQkX5Px5wXr2TffJEavuqMrKkfxCAHstX8EGOC9BWm/iL/o2kic7H+AL3ORnwVEzw
TUjmWqGQHdN+JTwbsOt098zQNC7J/8w4A+06vwHqHEha5djUKS72SddUDM8QMml4/xCF+R3X6klh
VeZqUmt+lCd6+Pg+MTYN0Jk3k2BrsMsQnvxo2Zbh7fvLgvuQ4mdQj4Z4XcqRWKcR086HgvecmPrs
RbPtp6xv8aw7QfbiiAVt/wNxgk1ZbCxgF7Uv5ixUO63htqpW6QXxANijlRIpBdtGTD8ZGhM5ZT5n
mJiYSwKTTGn4oAqco1vVNsM6Uqm92r1k1IyjfSOiLg3OEInKdIQZF1rjjRAaqNhIAUbkTfIYk9mM
10WQYfSV1oEsGRTSie60RAEzFdeYWljIU9yWsMyku0B2Ww2sjgCY2dh0rXWIP32m+U4MixWTBKYT
/2wOutAUzbk1M6vA8zmRRxjC8MmaFOeBsmJL6G3pcF2V8DMWVvc6WHKIHhzrfy8R5i2gqyH8QH66
BHmsDKkcEkx+9nQBdaZIBtONOhwO9dPgbL3mYzKrj2MzxNNVXb39pu5VQ0pujX1TuO/nx62SwXM9
SO1ksVRRQGKPgRMSIpVMKrzbpqmdQUhX+vC1EHXzYKN8o4iIIJLKONQJwAvQtmwJQ/qgSllX9lDV
9thDjsZYwy59FQSjYeK3FCdgAKo5K5gAQ+EthlhTRZdhbCLinDiz6Wvy5JalRfexLjt2+IBkFuK3
BZFUvmi/WMBIv5AbsohGiXrtXoQyNnl5OeOZkNReFcruf3mUtJVvxnNYjQPE92VYfNUwt/BF5jJU
5FrcEV/k0Ve5aWln+ryIPEtO5LRZ/Ag8dAcL7d5FMoT4dDROrealnYE85mHkPqqrsIH9m95AV3dI
pgORN3ns7iOAFjM7OApESsK8V6AfS2n31g1891Po7EWgkXYuUqOR4/KGu7Vd4pNmjFh4mdnVNFPf
n41vxQppfjPNqHbPPFoDg/sIGApCV/C5ikNT3VprefbgkXm/i6GVIi2OQRSOnGN2AMNc9NVuLrz7
90INSBpX/YpFMWrINPngUVnTpBcR6uO/6sPNEDaLEHB8sNIQCTXxERENcT+m4BwLsqwtoUfscAbO
A6LFcARZ8kxtL0U1PklbbPjMrSJ4TwZvjLY7qGbuYwvt5TZnKUVZ6cwgX66OvPHwJp/gbqDI97zV
xsGKAteYQhn9q+QICmNAPt3/nq/VYeCd6tbQ3/0bohX7B8r+F9jjT/auMMtdzw9bJ93of7SQ2Ptq
lsegN+UnL2OaWem4/TNjk1Tu32SGb/s987CHYgQRy4aKbmb2wynytL/qBGhPaVYdz6sMWwSOpELZ
1jqDvHAnPQr4NeomVY+G7YI7rsweurWQkK3JzY+yZY+jcRlC9I0wv/9ItEgRMbkEh3NhaQetL8Aq
9IQk45d7qVhPb/Y7XF66xJvL/3ZbPcn6czxZyiNwUJE6zZrXsTUqak7d/Bz6GBa6jcjfDMmZmBgg
SWqZlHn2tOBaKPZqyNl9Zv4UpFcnhjvXMCT4pUCyax0vFjYEDJz3a285T9MarttipLb/VHEATbeq
OPZayZs5PJvCGo1PxpJ4GCJcFB49v8AHdyexh1M8kVbcXgBGCl2V9BVV4Xm4bLcOTbF6jrpyDTZ9
OXjr6cy/yqVuoWsbyjvFOJzevwicvVFCf8kcQrhxBvPptRPXlx/M1/SqGg867rLZrToJDyWATqM5
DRfK7rGQ79gozwy3LbKTz7bX3iN3OsO02hnOGFTi3Lr58pznait7wncvfvit9Cjv7KNRXCi3Wy7l
zG942foLH5aQ2Ej10zZfrZPaBN0th8IrEnHtw2R9+99rq926gAiCiRDzj6D/RnpC+GKj9IV1Dooa
RkfGrrC9ti1EQt5nYfgA2LhZmPFw3BJRMNQMTh1L8Cqwph6abQCC+iiUAX5k8+3kP30hyiA9Kcyw
5+S3hpHlOJCv1gK44rYSyzl14ewly8SiCiKmAkmAfb9r2gXwMauU/7dBOXn+e1Yu/BnEKu7WhJpn
ZXOQ5FDj0BOQL5W2nE4uiehK4EUjBH1QkzhtAbcDWzojae2LPNUBM4QpOuX1OQJmUY+4EyOR4FyQ
nqSx10xOxiQj/EH5Hn4QIUFAhryxDWxQFgCgMK/P9ToxuFH/ZJ2FA99ArtwoD66yiK8LrdXuLv0a
WJS6wNVf1i46mby/LXyKTXCPHwp3t2pLsYhEO/e5L/oP+n/Z7E++J6PtGKhgF0cG+E4eBtavlcFC
zOCU2cQJZ+m9p/GtT+cqHhytMy76N5T4xsModcCfDYDm/w++0eIN4o+qs5CwqO0dDbG+AhzrhHd9
7MajPm759quY/wF0rX+EfnZnkJuWD7WcQMKvE/SUcDR4Hp0R/45TDKf/qGas3OEY39579LA4ETM6
+3RkDQqQSQH9DqpO2gHj9s184RNF5ss2yREoy4SSxefSpRD31+VKRECUJQWYnqH0e54hiqjyXy2W
Mu0iOGUFPnTufN7WrD/Xt+oOPrkpZq0pDJ/lOHq0OddNwe+4L9WmPYhMib5PnrR7RcSfIIKv91DC
j+4/6lxsfQTj+pDwzplliRhCnGrgAUL/bslV7hq9agGQjGB9mrvDRQ2F7JaKCyb6Io7MVMqdaYo9
NBGOp/PBHfwtMl7LDcE03yPElHoZ5BNcuzgSIMF9cs/XNwETRR1+fD1N9MoDWvCMgg4ax3GtAnmq
f0t65drqss8hOqBr09/0lFpUh+KNS3bStHS8OvbB1tC2kMXfUDZ2eqDwVMtCQWYL6G41KRa3apUA
jWqhSQikYZRQH55wK8uP9B9PfcWzHCGrcm6t0Nq852g4TOlmeJMYkfCcOEn85Fon1Sj19JQSmQKB
Agziz3wbWl72qP0kROfdVRcEWMfMN15doIJow454q6riHquCYg7GaiB8B45kDp0jkDvYUcu/qk9O
Ky0pGIOm7IMMA0j2lhFGGwDFZkudJciD7uAN5bJQCJJArFSk5nzbzVe5ezFnys5ZVCNHwzWT+f6J
6mu7RhG3XHTOyPrl+j5y6MEG3pmVt+jqxwRGAjUH4bJx/7CVPcui+ycGFC9i6F0EAu3hOavGDvgE
crOO+s1I+6ik1xfLGP6kYK1SixbXxC6Xw6MydeM7FWB2ENTaiWPRPLQ6bUmPb7/mx7FYNKWgYkPd
J27w7g6CDTwSjXIrR80rbMBpOMoBbwTzBfdsQ/XV88NK8zsFQrwpnb0B+0k9eF3EXOnNJ3QiUre4
vM9BeB0iwlibY58TlIJpTqKKS+xdF8gHN8hOteyDtHtLe3SBMsIajBsBZvPS3Nud7jFVRF+A+x1f
9dAgwDCh+y7app8fvD1Oeu/3N9boNahqwqyBY7jJxMdj8m5xmJwP2i/9tgV6o+3rCrgFIFuJgxoR
YO0T57NvnbI2cFcgjTCDgKJbY0FQeduXgPjQd/S3EI21K41iGPKVOmLRZhBUKCmyFFI/Y2W1xu0u
IhW/Kz+J1bk3qCpgu+lCS37Z7sZxLTXfpQS+SOoVFQoe2MHWr45RbPkv9yMa+QfZbhweQQoy3b8e
SVbfPlWin7lRKPw/1Kqg8J/4u8rUv5ZIfMXOJCoprEHqIN7Os2o/LuV74rNY94jIrWlwdqho16qs
WZD8mjZPsvd0Uqoi0xQRSF9La0FSvGh/40rnwXiMnQxxIRO1YWQtXOoNra5JN/AMSAKbSV/S0S29
x0xGrRhfAMYRoymBrZcmFlLTVbaFM9use+vDN6mbkqzTIfe+E6+zmY+PL+p3kFGb3dEO9zwIH0pD
5oCb2cNXZDWYUD9yQJ4BBlB2uJNl2gp6EtsbZJdz82YOL//+YdZc3ixhBuzlVAOh1vR8DBK4R4Px
vx8U6NSmZWIe3yEj6J7Svkoo1QznYE7n0a10QEUd1DpPlvlHyfCsZkSZtSXvbln8fZeiY//9QuHy
1FCTHfsdy+yq2G479HHFiKJzjz+49d0hiY4SwE6d9ecGvwV2IHQdXZvCn4JYgAqMUQOpfVqMks25
WvfCS1YVCB+ooeFmSZR3pqXkouSh+nYD5md97b+7RC6ufuz8q4uxe6NfXzYcEQYcue47hRDfUBE0
igo4wTTkoIB+PYN+yKr7BkBALZNqufp9QRFOxP4HyeFbn456DPh/w+YSz8HLxuPBEWPV/nZCmY50
MbE9DmvyTciftD4SKKB0447GQn6AX4xiNJOOXkPkOlHXM1KWdCh/bw4o4pCmBgsFXnAgmpPz2k8J
fDkVhT0KHUtGwBHs/n6h7Ryxwi1nHhorsqfYe72QlwLi8e8f2lP1oJwyufyTJ6M/J85Hh9tYrjb+
7r45Vszt1/9tq7EpkI5YMX3iEsl5yXOi7AZ/HCr9A4iM4RGB9KpxX0JNFIAlMzpz20AbW/YJnnLU
qf/bL440a6R+xq1a4RevLZnhcVaNQ08BPsQmkqoJCQEAfwm/kbDriDdjI5pQtrM8GmwfWcX7M28M
yxuaDBS1ewsP7MVoQLuOnXUlGW3bY5ABV7hDpq1W/0f7fvI9Uv1rxzbhkJ1orEZVezPSyx6H5agV
51QtMRD/2644d+rbRpZXmhpNQODIDLaYddB62fVi9LVPfIA1yxaWinZKrb3oUmrD8PmyeMwhjH98
a5V/lIyMq0+m3M6r2XQ8hMpWqTJxndnrTXkzIzuE1Giwq8aGBqxQZVd3Kr5fR8OIp/de2+McSdPp
mDHVJ/SgbMSt6ExkUhS7FUzwavQnCtNn0zbZcug21q8pn+YxRpGIMTVFoUVuB0wUG/JJlJ4ikKYX
5ocoSBBtt8+Tf0eA485Qscri/Ta54gqVvPjPezu4/+Lw8D4bAzBo2JC9e4TiVA/7aWAzE5b9Ys+5
FNzhi4myZlSyUJB2/on/1ceIdhJKgCNtdZZPY4hpRln32ZH621kX+ty6yehzXHnoy0MicN0gPQby
s3u3vbKsTyZsaOpkoPE4NTk99ZxXlR4ah/2W7eHf79/mHlNOnOyI/MGmGwJSVqAA9zlo8Wz0ewXI
BNRAwbnbCjoKBu1PwTdFiuTx2npHGNPvaAkn1gOQL/+fPQeHe0QlQaJ8Fx8u9C92B5kZtixjcS+b
yfMIPj5ZAODflcJuepOhXkovx1pFA20a5hHju9gNqeEjqIeGdThcr/lVYW36LAsvDzfk67sfYLy5
6duUQrVupSE+d4+6pf+LV0HHawP+XuxYsXjw6cQjMq7CnsU1t3fukl65oLL7tHioc/jdQmqEpVgl
AajP/cBpp5pmxcnrGJ4W2O4MwDke+4g86qmEjBbqJ+i6Xq/ks1VvpKGcOY+m2NkI824RlB7JydL/
PoLyPCkdjITy+4AbHPDQpK0QsDCXa4SCs1QgrmxTco9dXeL/50Ma0mYHKsa4Kldxm5moPHH6RfNy
BKp5qw/6m0aWsehJ8nVjiRoddXGz1PtqJIfgrTcaXywzUknoi0DtmkikwYUNR3NehOe8mg2bJOtO
EqSYULyp6orFLz/RLgv96dICqOLwfqTjQD5uUyHPj3Z8WWWlaP0e2ckEIhE6OckFsCqiM9ofg2i5
gKxQ5/2y1uSfJyzTxA53PrzT5oI3cCuZJQRRiCLiToVgdRFQ+5d57kqR4srQhR7w6r79aAhaYSBS
aUvsQ8gtdwG7w0EtJ/SrEvf8YAM9hWkcfC8euZB4EJr2g5x5e23qnbya6Gs4ZbcqnfIG9C4ppg0Y
TFh/0v+lPsG7HShKgRHeSlV1jAj88qmCZPru+u2QiB2IqgKuR/KvCZScRRdGk0MLYzAhqpu2xRon
W3oJgIuoxuc3PY7XHfZlDTOD5wzjm5/ZKge+TclG0cvHKeAs5FnEnZUYKFnmWgnXlK5Mm0tNFk8N
RWYU8OuoWASR2Viok3REuqxS7ramX0aiceVqZ692WzKHLvDNWT2l0DisZIr/JsMrxS11/L/8SE9O
An3SXc6pQWH+Cjgk2dHB8wlS2y3tV/TZOtoIL3S1pbQsBWD6HpiOl4SVxkWVlzby/IJCN5AWFPg0
IX4aRKAVr6Qt8S9yZfXmqUzE7gCd0fNdxa/zk+t28dBoDBVU0uCGfYIj552wGU5VM+OCJQojZh7G
J+IVtm/iEQL/ocKkYd2PG/3iO/toz1yH3XdN9mi0psCHA+5QxGzl8g3AeMR11ZtskIl+yq1178OG
20EI1oHogAN476lvEe4ZPFTeg8SEVnOBoUsM6xDYiZFJp8fhjdO+Vro0QBd8bOoQnmENnxnQhusj
HvKvBJcQOF2AubvFhs6oIG0Iy7mO9c3zS903c3ml5Iz5XhVCpffiAl1WasL2cZKUl73jzL0yb7bo
sns9p4OMxz61bAYyzRnXbQAH3pb7MfyIwWSjfWhDREChY+MGhLFzvPjPjc1C1Yxu5dqNUuVNjBfd
DZVmE+jxs4hprO0ZjMRR8uJRe8puKR4JdjTF8IukCwFq1vgjDpUxXLyts81Y7f1ErOSIWaZBW/02
bv9Lcrkt76w7LSrX/1spsqV7b4+8F9M77E4YO0ehXOva1s2fu1Lcf1JOZkpNk+wEL2VgW/WVk/i/
6i88CWSxANZBDmkSnQT06JfQN6nDVCz9SW8uXEoD1daqVYxQ7Bbe7rC6Qf1WzIWnVjtbm8Llibu+
9FxvHwqzLnKmI6TeBE+pjRdrFh8YNJp3l9iLNHPzXg8OaJwsT9WonurmAtG39PCdzuuIbyPlCTie
bCswi0C43zm+sKdfRFfEOh4dhnokhwx4cCPrwnJq/2OPJOpT3bvFYwQn1Bq+7L9Mj4Gztqg+DIbt
dnhOtCbH1SddYXS/x4JzzLPAB5mCddpR1WoYrfPOctXPBZXSI6ct857lb5/A3wtaiW4/n4MkmVWf
CD/HACzFsd5vvhhLQUpkxIT2HRF7p+NMFRGvvpe8CoUfqdbaiwiDD3g8wvvFAi2TmSkvZdOd50rM
NVeRvXRL1+bTiBp6eHB0cQMcnf/+EAgleTzijrgVBCLhSJkB1BXJhLUf3D02bZUCIj5xcBf6GZD6
Y+EL+EK52shWgCGnRZC0Q+5kG5e8IyxSpoCkyo8zGoeT0tlZdQlneeNriofaDenVu1FnT6+v95PK
X9uua5W39V5yyJxSljbuhLBbm1LwhrjC0eipA1/xHYYFrDBE4QBIVbHyZfLjH1t/ZPEL9L9sWd3g
KGkMkjpesxdsrIGPE+7vdxsT5auY7T1LBuTEQ183JjnDkyLtwoQ0NJ0wdqTWZFHDbcGd1FnXXkID
pZ1co3x9nxnzyMxP7Tm9G+l3Nmb7xsMv0rxKjsIDhlwVMgazJrjW8+DzfEtbJI2AAQrNfNELrikW
jFF9YyJCXsRR1g1RUYPWcE8UuM8NNOF3VggnBzCeKpRQEISfKA7YwkiNGhfLNpgAZcllrh7vlP2s
IxZu1cHDMMyzmM6BR8FHBVg14OvUA6t+VMxiwEx7666qpgW6k9ME3aq0IYWvb/MbzPTRJWkRf7uS
Er8dTCgLcyUZ+5jmI3vrPW84jxztvA7o0WoWp9ByxfRsYx5bKJsD/XQ/jfpG67Pa3+z7H7B3hwul
6acmV8rMMvqwMy/bx/7f1vp0PfMqceAWCLAwOo9Xb4Ts3tMoSWEwGMiNAeHMY0kh4EHBIh+3Zspm
CHQcZCIgZnpiSkduDRNtO6TSBgp/x6DE+hLvuDnfp2CqPJbW5H9GKqEl+Jj0MKf8QimeN9r+v7pe
eFwsLk3GTzZ4lXtmIxUeZYMV5AkHvxD7xrV1kjBXmnpMXwvUNG+su6+Dp6uK5TjvzkW22c8QdLgO
fuwj0tY+DGKA3OjVtHnEwLJKDBRxoBdepLQvr7MWWrUg3hCTar37oAcHTje/NGrNPNv7rNX8vKud
C1vFJG7VDKPQHnoLw1jmeLCn6713hwRNSXmbeQ1jPFC+PqUKPzi1zrtLqXM+Ma7MULJusjDC7dMp
qAimBkw5zWOv/Y5lLVra5WNLpiwJstscQWN/RU1GtfEIIp76A9qyM/W6fBLcVw0UXh+I0AcTRkXf
CzC3qcyhFwrjoNg37X9y/nXHDj3VMkjUWBCi8FjkEMotFD0LpMcdyPvv13K/m8broRpEY0gpRSYU
IOYeFM0l4UPpKW4PSYaRpHoURqcmzko1ZWITyljFnXbnwY1mM1pIYNsGy62lFUoRsuIOcERJQx3k
tX7+DDACbAYASX9YpJHe9rCEA4K5ePwCdqkJrnoFsOgOvZfTRFWCPMSgaWt/6yFD829bf9QA1tpU
fFYu3z0BH+srAuJ/QgkLm/eLQWSemkzboEIJgoXeiBSMFDmRagsd5tiTsII82i1zT6PGC3qdTdAe
fItdZJyuLy5OoNbtxX0AJqhudpVUuvLFCU/y4j3sMCo9IGwSd2LGql1Lgx+6eXW/Myzgnnc9h25g
ZQ4SSPBWKWtbnJZlFBLGSs3cZJT9GMgIm+D5m9QZmtySGtzWzwPm8nAHOvF4ktM5+PL59wjGGo4S
E/9vSETTSfPZ0Sneed02ZNulsGBW8Umbfsh5aPqevzWdFDdW5xItP4cA+v0OnS7VjWUb0/sDNSK8
S/+WQ4Nf2Z6ks0VU6fHMEFygCwY3irwg4G6X+nkIBh7gI3uW5AR80FTb3PO8zkMIeq0kfy2QJt/m
kxJge9c2RngjobF0OsBgy3ZxeEygW+hYuVCEp2Ik+E5h+jkni7z3lDnD1vICrmKAuRLyD+xFKAuP
W2+UKgCZXvy6c3WvMLrejsIi2JJSOKdJ5erEmw0U5/He+Ix5NU0BP3zydUdzpxhlT0P9H6Sc0+fs
E43GEJNIZ9aqn7hUPajZSTt79G+GTYRzQ6dM4xr7PUPckedR4l5AhkP9yPm4V8Ulcmq+GUI1jclj
emRPsUZ+oM4tzAWLAMvewfx+bUYe5JbRxs7HEUlFQYmLOXK43teVZ5N6OgWSdgWRnrNTKP8uvVJ7
RTsdEnyUoNVUG60piFTakHM1WuIfCJ3eKifwfQlxFAiHwC8vhg49uxacarWexI6ojyyQxdJ7PJSl
7lbMcqdk1tGxWQ5KMSxqJSsXD9Jq06ilnKG8v7qyn0UX8b3WuxD2f4ZZQRMhSu7DEi42HI3lBB2t
LFkcFGkhcDf2kVRrTih0RKYlwmmiVM1Zd/htAHRmOBr1ZPMZay+/rUn0EBfGfK+M/i0a7w1v0JJI
/NsVKKuQBCDtjkMVccLusOSQtH59XgGQIz5zpRU5cbhIKdc/xu6Ks4bhoKnhR5flgYyv12209YUL
kamIRae4Mz+2LVdkMWcTB9fIE5yMIhTaOZ6+pt1cW6Li0MJBqUU3Y97TilOSG1A7e0TTau2m76zl
80b9egbtLXI27goL2DAr4oEGBRuBa0x/IuTYvORh3bBrV5oLTz4pF12OFjhASzI2gIXgZb46JwG+
mFFwdWiKRZvABWs0AeTeXNd1vYEXKAcTAvyiY3LHNG2W9c4KpD3NCjWNbAufUXtEDN7cBlVb2vhS
8g/3a37O5N/4sJ75vswp+PRKYPDyRfIs64TBgDWH5JPq2lAJNZd6GG+pGdZYPfb+aWxxIWjtUrgt
Xd69TSyhPA5CKMlTgpFbrDRf27q6l5eWX1p0fKKVPwyHqJHtSzj11MzRE3MRyaCIuJJL3aFCvMk/
drorCMaX4rR+wi0YINxq8O0YY/A7+E7jvnCjdwLTox31m3vfRQrUO8nR9U8Kjs7n/IGi4y03k0NI
xQ9tWKJN85xgTKygjdv2vaNMy8jLd7Ysmxz1ErqTQQ6VJ+euB2BBG9HznNBVIPjhLVJRE2CN7NCw
K0k/s9Rc5HaRwXFJRDkHgkLdIDq9PfciNOW42je/yUR5wLupSkBoXcp5E9HjeyQkjJNdNARaFCx2
UF6i9y4ahMfLGlYN1WOIaVx1Lo7ahhIZGRUDId3JbRb3Mcihgj7OjRFz3H9qevngi8pSz9xNjiS6
xtHd8O7/YRWjp70Jx/9iTVX7Vres30Jqdd+3CDtKjyeSpgfDhZdSAP8VK9W6Ru9gcRztQNDyHrdi
rj3cHY0eO+k98wEgWqn2CuDKfITu8ifhPWspLdOLIqUbe3CL68NwZ7TXzFkNKvt4UAjEELkUEIVs
sFjVFoGmvPe5QD7Y5iDntYNevnUfWgtdOpRaiMUMlYZFADUiIZmVZblTgL7RIlz58zCIih2NgsAj
qI8kW11GXMxbI2eGG44D9jZw70o+nJRd4ce7ppUeeBIeDYHJ6MqA3HWXG8MuWS6FL7o2fX3YM3KL
bIFnKXdmQFb9HMzUMk9evD81qtN9gm1cA68QrZeVUY6QZC+olZyr+Kawu6u2dRJkZDF6hUeNpM5+
BPv2r6MpWZuevQB85pyrPMl4yFEUo4MnaB3p8QpM0hxbgt7mo95FFDikZePGO7dVer4UCpTzZaow
EQMyl3gwzPFXBY4LM/cPDDgQmcI/VInkUwCGy6kjrRf5fnM5pSpHUH6gxyuaBDsfDBq3UvMLcLIc
jUBvnAVCBZQ+AZrX3YG7EDHSCNqae6jDgLc8XfMzVzpACxc/7ZJ4Kf0ejuijyPybjBq622DD8Jba
GxjfyByTBf3grfVIqkdpvJTGo8GkGVSo6u91H4rjJdbqQhtCwqzJObAk/POGHr15P+fswscnr4sg
61+UOAciOJD78bhMn1+tRLZgcCCgCJXMbNCIbPC/xHQCvaSmsjSg6RNFQoFw3WGwYveSuuuP0lT1
SpTit9+xRpE7ULf68olGWd1830DRsdN8AE2YSdQFgsRjSWvSuAnhvc7GgbLNSjC5jq+TDPYSBef3
CtJUNpz99nr60FFQSMpQzIlwuIWyuvNGU0xkQoTaVhKsXjkLbxw466IKHib4tME9iAZf/NlyjQve
nQZSeOyVk5Ut9FzChnhDjcXnJuWnkf0bNStKQgQUXBGrpJ5xOfvSDOqUuQwfUGu8fI2LOSi29SQl
egtn/Itb8obI2XJAD9VER30Zu4chs0Zxbkf9r8doSP8zLdoMDBJFRYAZSSbkWwY7zYh4RFXvKFjq
FUYv4sFXZgm1XxH9sEXdB4F5blrpRkv6YtGhOZ5aORtMf8O5AIyXaUCwwWurFOLxMSzhq205N911
vjZlbS7N+hHBgK+IiuXhC0O7TOgcTVAeGNFQMaGu9D6Wswep1Ph8/N+CEAw1pK7toIuUnvD6zIlT
hhqZz0cd/W/XpcyOwQvlywPzQDVcsIfVujuKen8CLi09r/hV2H92a19xB6z4tPS1j9DjHnUImFfS
K1G3EKHevLOs5DN5Ea7DOFhX3nwKaw9hk09FUSGj/jg3yLvD5INQ96HFReehl/m0S4tAVfa8VVpk
6hMc1QuG7bz/Jk+xyfbINq5PBWSKd8mseH52ORCPTdWBe5wpsqXcA1NXJDRc8o0SKzOPlJ4unIvK
lHEkHNCqNIHjFdgYtyl1lHpU1tuoeOU1SFFKPzLOp/+KKBcw8lbsp656hAtxqoa/8CgU28fKJS+M
jfAuitfrltzqYJUxOBmRinAgUr6l/qv9sVScSFhqixwz6hAd9VVbTxwR5ZY57HcoGKFQSY6ijZKw
UHkbmgjrlSQ4EG8ZS5apwrti5dSk0iJj2GWuW7Cd+XP4cno6W2VRVm1wFiFMmNXWvt6abe4JVzCd
PImOuF8W8UoZiJsaDxmg0gZyDiYdUiqkYAoW9yv/+nJN36jlfn4aUUJ3JGL1xsT3qXhwDrkTqIf7
qmbID1zKoBJiBjuoWJtVuUiaHx/4sDnq9i1E0rdfyrZyfqR7ci84xdkVJ3t3q3VLyRlv+PD3XfvB
PXTZliOWObXXJla2hk4r2sSWPNFcwu6+wpL50wig69XeqVn7MRtvO2o1/xBVj3aPn6iEKpvkkgN/
2vycuH++zfqBdc9vg1DIDadEn/d6cVMdpnlKyCQH/le+Wwf/Z3nwbd9NblZY4mSzu1DH3zlXL1OD
xxuJIIEj5joumLsjGpMPzHv+A9g6Zru+NuQiaQJkcgTAYg9ajPTcchG4iz1u7inP2xkNQzH0cFLg
UsWnaZAbkktQiiwDFrGOYM5NZsYRndUardsYLETLx7bPlpo+qLwSpQ8EI0vKmNXvyWnbUKbqX1En
9kLUiQDL3nwbMAar3fa4UcbXsJ39rLkX9Fb/2YBkxcDMizEiHfTSVFisq4HcKUq4o7ed0XgNKvNk
bl/Hkq8rUsf8M8BITDyI+aigfk2cWsYK8FPT35Mujcf7vRTGdosLMFJ6U4jNip5Bzy1qpnh+kgQI
MDvLyljaIqrHN3RQMHUmOcDKYa4LQxFGz2GBeq8WMpoloBYUoS+vi++5RYqhceINC9hgZI1Btflr
6KYdUPitazj/TgROJqMY3xG1CYCO0sgVXZjM+1UBj6856coY6knAHEJ7yey42SWh4Jv+zPtJwspN
8iIqxWr8RXT1GjfFUmm3xflxSFVCJv10RhGdGWrj2CRG+X1yDHLMtWOejl7T0BR1SB/9Kt2LcUXx
yV3KbP3un2PiTuBMyhdQArTkoIvYUzEe+4CgS9mpGijy7UacOtCWRF1pMpQBuh8xcFVRZ9gZMb9w
NvOhuyJYUl3w/a8TMlCucOe7g3/d0ip0Q17Y5qjCP1Jew/Vx/tOzDH8URUB0kty1IjBaBSTE8QWx
H6dHN01IMulWjZaz32xUnttOs5P9qFo77w6AXFcfUOMDPIMb3y90lvKLyB/l5+gSM/VeinxUpWRq
HeF2aiginOE1MRbacPobW+hc73YLxNwCMAxTIjUf+rbLas+WYRM7cjlYXseZvMlYn73epfMHF3lo
XRMUj4FovBx2vs2p+Cb2LPTFYHKmYTlKcDPfbs85GDdsXpESYzXVAgUD6nJmykbzEsmqHDg/IKv1
omazDSW2HKCnN5QQ2B0ecLJUdV6nIlIAPCn/2iAS8oVIHYXp7NLoA4qYl6B9vR+PhTPTuTZnXN6p
QcFBo7g8LjvAHP+gjht0napERZAwNkV3fKWKfldkwZyydBVX+0jdg7imOY4zv2H66z8aUrTd69Gc
xEA4xRkbFDQxQEfzL0ICpYK/STE6w8QNxFAjzubUv7cmCOnRB2TE40SHBK/uXEtfLqNxq5PxVRwk
2BTu7Jo53TdbWOxmT5BVqPbyeU93oVq413m5fNiyYL50ZZgZvYI3exop4iQ+fDMlgiaEkAWUvwh8
n2NIDn5158EtROXEstqkoeXQPXu0gR1jKZt7YNJx1TqKgdSvHJjfpvRxyuQe0ZM1Lkfynn0iVMSr
6HNDIu+8PUM8pdd8ezRwJB8crH3JG8kg2D1qY9lyB+R+asckkFUlae7Cct9r8jhQ2NYJzHySPWs3
Gylkoe90eCY2k9mlWKce2+arhdsIPjAU4IVSRqvnJO3JHSb5ibejXjSRHwnnukRpHbvSR17leII0
uUbKpTOYxzGfJPkdJB3r462Wv8bbmZtZ/+F6FCq7Z37G0AaPIHNjh9IurZDWZ2ZQJkGhwrk593y7
SdwMFQDqJf1ACOfFBZHhTjLS8Xro7ZjuxA1K+GvFB4Uwmkpql856zlrhAPxk0KhuC31CCdaW9AzB
Q9YhGKoPUb4A4cjCPqkLz0zd5KKFkORzMr7lt+SIm1G7iyS62QKtkLLeuVNJuOFGVDDlXA63v+F9
ubeRzqvFDn5Y4MNSCuFRhAEU/zYj+BuGQqjIhCMWt72uXyfOSeGB9cXlShEWICu0TP77MQ5/Eb8M
y3e8szDXqUBthFCr2t4PqZ7goZl2fdBJvT8o+tHZmFNdoNG1dN+0l5C8Td5//NyxzKydHd+w64cH
wSXBcxg41ZnILuz8V34FDoVs3Yj7zj1sctRn4xN9ZLC/UUmngJf80oMaoVwO1CrHWG+g22SITZC4
FSV8+tzcNJi2pKhQroXzS3hdg9UYgK5ZeHNGw395cvQJxXge7a1STD+Nn6qNhKwOC8hrET+/gn+Q
7E8lyHKHRAEgxemgAqmmw1BkKTQA5neU9+3RqZ4JiDphB4Eew/bOfiogqJGg+QM5IRkpZqddV3Qg
TXqZAS+J41cOAh/S/DB2Bg4tJKr4tuwNnE/I0XD8KztICZwQ8xxBeO1PLOMnIILm7LBDmQryiRYA
57A2xOZnUjxKwmE+f0gzWSAAC1y5hNmZs0la2J4xpBmP0W6zCZjmrjZB0DGW3VO9imomluXJSZKb
rdTBG1vIhDG6pevfqGOVxRAMWQjBF7mQ2WD+VYG4RmUnaLxyMNd1QuLyc7BjBRy2+ew9PcXJfQp7
D2INY9bPlNd4QtjWEndhBMNzNMK1Gin2LFRaoEU/DuZf5lwjxyDJIrl/1Rxx7ARYDLglFiqEJgLW
+A7nrNKmhHhi52uoFkWOg8CLPzSXhscZ6seWZtm9vZnleMeBlp6J/uCqLCeEg1bTAKCgCHPcqmgS
dYLCsMBpUi1fjLkRFSK8P2XD1jxEKpAK6T+RMJjMbROEcFlPHooEkDs6y552fpydDgvLaQglmvSS
wCPOqrPs5JBLviUOt7Kvs7Y5gAMHXBkmqVEvRz/I7tzD4Tc90XtS2/SF2Cek26Scc8tfvGtPJYmj
AMINvKg+P4O6rEaIdneTlmtX4y1cmMwhwZIf5uFh9hHRON3WsOFE4v+3pSv7BszQUPLq9UyDcVas
EmCTUWZuKo7bMAxyMreWx7k269aEdvQnkJ+BK2bx0Odp1qVvNWabnV9HqkE+dh1Sl5sWSW2KLehq
F6vYTZrOnDfU1vjGDGtfIyrA6c7sbx0Ek4eKT1S67xyFHVwmZnI29I3AShh0RUU7HPzYun772GAn
GS52qLFT6hhPV3uK7JtdT4T4Dsu2wcqHowQewpYuYta5enhab30NY740CCFExL+3NtIy0QRGLr7G
g/D7cC6R84wAHPJtFBq+lFQvNHpffsgXHpR3HP+uybWLlkC2pM5m+SEgCCxWjmLzkkAV+tG2PsRG
sJZkZE5F9NhopArGqscsi4ELRHy8fjVRLaNOz5ROsZpZycJV4b3NS9ttcbPMMrpzxCZZQIP4JINb
F/Nj0ykuW+MaJl/h3IZ/Ev53FRDodl0NMUFXk34Xa/mjtlqHQNnG3ARCqirsMq+Z2j9HXnNThJ9s
h0eDGlW48Y14d5KHbY4jsKCHpJccqoCtNPmaj1s954Fq0mr73R2vYUGQaAZMRDLEfYW3unOspxSo
YZ8H4Bvk3VrCIlD6aRLPKEH9E+DcrG5MTxZr7zAPeyC46hvXytpNxvKOePuf8DGfs1kBlec8KKV/
yQDZA95E+8tAam3LWThBJkOQ/RQUANRU1l3KFGe2e82C3Tzx/hVWBRt24BBV7e4u+4vSw6JVuDu9
si7StLmmfXFWE5CVM27EiB8NFBEOYsdrGxaDGNZCpyK6NRIDX8zDTx2TbaBXYIZ7+4/zNp0heOAs
ejgDCgcFIpFjY/U+km6Aihnaqb17V06wQs9C9FiUqpPvPw03xe+/q/Ed0tJfB9O13ukudDtDFMZZ
F8Z/yhADgI/OSKCYFZ1DNEzlAkps2ZhkltITM5L8sQrGsFdBOCDvdXGFApyoU+rvNeUEuXRb09DN
Z0Cx7+yVSEg9tUs6vwkzX6nGbyIZnQF4OVFUNMa6iB3mXurjlrAyViSFb8cmpGe/6lMJftXzYKXO
ajvaES7DfVvJbLv6LmRvGpL0gD3GhO+PCqtJvRRjX9EI0oIQqKWNBJHst7Qb96dW1gi3q/ZdZid7
BdIWL1Foh49tZRcvjLVSBN8F5msBVYYMYLtatsdhm9idUtqi7ydVpvgOaAAiy/6I/9AZ6a/LfOh1
Bqzw9c2Px2k2KLOkWRnHlYc0v+d6N6vOJs0WekP53C+8dCxHDt86ORncJfE9weJvPo+FmDTzsK6E
9RX4SIEW9zrqBtSeCg3D5LFLthychwd+2MHpsVYEET9EAn8thAGOCXIFwyJgZUX4QyJhcrlSHS1g
rk6jqCOvit+hliurxcny+9fYaloedt91bsRnICzhAAOSyPUz1uqumwkH0RKcJhDLgwr3xcg1PioH
fvhlyo31xFkcKCDHAGoDfpmTZNyL8reDNAFBTHmN3aT7Mv+9R2s3/y1rRn7SajPXu6z7+HMtZAYL
pRzY5520m5g5OK0q1Vc5IqhIKByzuP3I+OEU/4zz7mrc+scnjiNYpnc/xVTo7MjSvs+TTQjYeEf1
OcMwm0/rHwcca6LM8op9085Y1OkhybxIhwKMqdhSeaX+Iza3C98wUO7QZOJFVk5BHG5fQpTCKLLP
fGVT++yhp9oeGEfd6qMD3aXeDZ667GSrnAcX7f3Z/If0LeDiU/C85YwjUQWvzkNCcEGHHEr3U4UE
veK1Y75p81keksG4RG1HHJkkiY1EDiIXsfVlqsJeJrCHX5lMZBCs1/LhkgOPH0WLQIstzBdp62/z
5r1CwW3tVit4trfI7ekVjrMpaw4CC+6oXKzcPOTYD8SFD/htRLbfvmzCindzr+wPqKJSTSaoa7To
jvqZrbvKRxKWkZYgnSBfASMxYPBIURtoSQZX1x97lq4fu1pgVJRHTAV+GNAKbfrJMajao8YDkR6Q
LYotqwGGtp5HmTWffVdfQs9Npw8z9IgEKp8D/2iO/jrWs9+qrODq8x/FPVA7KB5D8rD6Nxdx7ypP
X+vdbTo+p3QdHqNRVs8MjmmDC1pdotBXQgNIuHwY1Na1EoNQagrrwnNGFn7DFdmUfpFEyg8sfcNn
+7TjRQBH3O9CYNMZjY/jexsoU7z+5eQI/jzQndMEhqaD9/olSwAcGTlIP6SNzQcHx5T/C6YYurS6
bIKmHU5KpuzwipTAvC60Xg+yVJ7EwhmldibW6JG0mvhdsRbvQcVcSONMYv9pUTfM3BKjTCF5NkRH
hJecq211p7SmhnGywZPVPK81LdAGao94GdGd96JMRgyoOz05ny8lQRZrUojO6R+Kr1ssqosGTRbf
7Khi7AVQFFwNV9l9jdfwZzTtAAZobcfFuZdmXKIXtLLubX0C9mts1cLD/CCnrzUfNRyWzsD+cVK9
Bl4DpkNR5u5O6wl5InHKoN1zw3f86z5mP71f5/27cZFXeX1H3cG2vQ6Vc/bEq6MGvCNV1nx8/cjp
ScocB46a3Le0DbZ/Lqfw/q4WgcILYj1gfULaYSfoHnmCG8hu11IDsL1/050fZ6KQbi66t/l/acqW
TFoJs3+nyQwfNk6pY7YBzTqkSHWZmMkrkbIs4GmRaVh0b0unVJiuI7J/yDS20S08vOzyS3fjH//Q
UxdRwhN7qQc/IYBWf5DxlQrFzNJ6xqsV5/embar7j5l6uTUFymxtcGjUYYLWFN/NnpD6NTMIo6h1
6HeZrXdh4FUTcgI1otJ8M7oCiVMbihYCuYxUK7GkYU38h1UNCZG9VLeZKmZ5sxBnldXYNSqDzobH
txrbZeZBrebJFev5033DidJ1IhsUP8mQEUnGysnwbGTgJu7OJ8uGfqf573XvddmwiEpPHqq2T9bg
HNpT2RKbxSWlQFafxjZhLKv3XfPc+I3enKaxh6skLmIpv+W6sbOXz8RRtaq5TfJDFSokMJwGOUuE
iOoCoQ/FYYPTQIgw2+gA527lWNJblUozslS67pNP+zuY11veW3n1DvvWJQ/hdsMc9ksRilIOId1k
uyH96MrG+8mTyqcPeaS0vlNskeLpgJpyXkmyT+FTYnKqA41gH5dudka2zqESZufRLqJKYJ4UbQlT
rlDwcSl5GV1Xhf0aoh6yg9uVW4biTWCrevnj4vKCCabHOGshSu8Gnc0tLbwoetAeen6gqCIjDqy9
E7oVdo1+okIO/jGvhwsQyjWRdb+4yc7BXDjqsckvA/v4zxhJL9NN8i/9afZ97W3oxzrBWFQ9ntHV
itwrC7SEuqBBsrjyONIZREUYyB8DcCSPhiju0+I6ZAM+WDYHzKT9EXeTjl8OGzHqE0122+WH/qhy
o1KYsrRzhnPY0/tAHvpwPzgmo55F9lhtT0+/nI8csLtvWJIM0XgJsOZPpDOUrLzcUIp4QdkUVwKV
rwxGQ1MW8U37wSyJFU8/eRpDowpYpiPjTkzs8yF+xIHB72PSz7FcZMMm4dRU3BBGexNA2n6VDQop
2Vhwq+7pK1Z6mH87XctSpY2TCYuYddwdY5eK/POO4wt+Wnf1KOga3Z45Sx9b8PhEZ74dw5uO3/K0
+bZ4RT9MVSjxmqKcKaNwriL1gny5CuC9kHLLYGCP1aUHQWXsSSl0wPxliimsGNn2H4meXiMtNn82
LXDAt/zkiU8bWWteGaPCWNU6aNwheBZ68Hp966R+3qDkHtMMnMqp3bTqSoVZtnOId0X+nJeTiU6W
0qC2tZZMrRBMM3fzuFSfu1ktIVh8dCVLCIDbHuNMU7KpXG2C6GDSjdnvEvCZnAWPvYeKYnEOftJE
X6IB2mMKpbIENyAy60r3G+NcAqHCyuwWoAMrrAV/iwNcTwjWCdKHjDruBxPYAdZzC99n53hjw5h9
ES16VDay8goiNp0rVfCUrnQQXP0Q+Mn80Gx97r1itvdyYmGhFcL3ZachOrszCX1Spx7PjPNXscB8
5T9p17t9AoreX0HNzu2a06X6PYAwwxDTDcz2LJUX5T0e/qyJJt8pXO/j6523yb4IBHa/Cqzw7wQ0
GNUGY2S77C2dtTkfgeBzk8FOIpYVkndSDq1eGJdWLe5WQEUK3givTw3WthV9xIWRzWk0HsUHyr8S
ydoWgMiSLOLjDpFmk6a55lxStj+AMBmx3dR2q4aE/xHkUimD1PcDLJLPPPO+AW3C0PQaOYlXt6+C
YJ+QLSTwI+jIfGFF+8hmmUsaK/+Fe9jh5qC6/m2WOq8jfGtP4gtrxw63puq7yqkb7hTIzQCINjcV
QmlXIZJo5F9oPcpWvMJquTblMsCwHV1NJwgyYDPQko+Ldh6RoDzK6KJfLW1J6zFV7WhYJcJA2p+L
BKi/Kj02z6pseTzO12Imo8Vp6fmTTHkigO551zVAN0KIb+EmN49G7A1O9bO3FRh3enWN0cF0O0jg
gnhUuelQFqaR98YwkuxzjQvWgUzAE3Xv3yOqczuVFU/g2TSBrBhBfgAs6TW6XwJrx+iDugCcJXzN
JEacSNlBcE+FRcjXK18p06OQ88Isb6qI8s3/Keo0+N1n0n2/ahBUuQ1jlt+GpUIHdpwvpVMsRIG8
yJ/6x5EPKafNacqUnMF/oeoBeO5/VwivIaTI4vx146skjTqmsGX/5vh+Xm5ViySrxKN6BWnmVt5/
bf5uPwl3jPyEyxBH5i7EsMAJHfGgLglVO5uJ3qxocWlpyAYySaCBKofXRhTs4C1diWRuvDJRSKiP
CUNp+p+nCK3Fn5LRyGyP6Y3nhyEcz1XGRa43Cll7vb5p9yJXP80zkRdRhwmu+8904CNW/KbngVjA
l36U9f4NCB/v3N08dZF/zS9OpkAww4wA9qGLOamIIiY987zNKsbo6HiH8r3DTEHk/C8reACJoZID
zhfOV8bHEOFocmZE4JO5NfGmJFBlCoCSQ3vp4D+BZSVq3eqo83ow/cfuaReUketyEiIfx9+fdw1p
QTxp887S4uybwC7EI8MfXLovVfzIJ/KH5jseP+c4sjrNDP5jxQcGytuyHamBE8IKdOpMpGYmjT/p
/Y9sHsj187b51QmtcfY/HPG2mb5aCFkDkyu2CKZY47BfEuKSLNZvK/rCGDZ78wOAak2UNa1Wiv8h
qUb0vpTQtaZjNhhEcJdOJ7vcv5N3pMGBQtaEKLEwT+h8lGKKrQH22gqMClK7rDf21xFygjZJk8SC
uuBZaF5W+HiirTxC8nMYWqO6dZglcsJoGKxvQ9CJZ1UXDomNC4Yc9BgPYygcs+MioYrMznnKNOcA
0B9MvKhzpoUtB/zLZVddnMSkfDIH5sB6DJBhLLZCrDivLJDlNZEFBa9cvQ5CuN4oeld8PROq9+Sz
62QmOkossZ1MlbvvhcUndJgYMzAdft4lHWl4yKnuyuV1BPWyPEnfLciNAfpJR+R8vntM4xcNmL6m
WV94Ovi3yAgTfgBBq62BK1pL/SbnMaYq23ZYsGPqUfF15LwYXNo+K0uyMI5MR9XNXREHYlfziO0X
R9o10k1jnm+rhWixvpi2KlbaDVF3v4eCINehLjJZzZv7VxzCj7QBLtSPjQX9lAaxNf845iuiCoL7
XEnALTd0rkij6R4q1cXU0CZp33XsORw7s30sLSG2zNXolgPiaegYHObFTYLjA0Yh5T0wLIHMmWgj
c4Kbz6JueO3R0ejgbN0xyp1DE7NFWyHCiv2g5v2aN4hDcCNWiGM+hUVpXH9kQl+0dEmOBbIZap8W
j7YjDUMIKi9ubrGh0aEo6xPlJmPsN8fa5Zq/8pMtk3JSvD/KoXQ7WF4h9scJR9rWfWd+yuuEBpqr
3yEMTSWuF7+vSdbDl53Sf1aQEmGl0HAxBh9rGxpcmz13KIKYmUdRlxmzmfurNLz6rbcTMGPFW/B3
UHzGPEQA3Sg3hUgjKdpwNCNxRJTzznMrMngNwZW1lt7DpeDiobdjcdPcHerbjfBVGllZdx4b4kvZ
JLlgd8FSvPWlJx110ZuJsC1PvCSq1UNUATUPMJqLe5/zymHNmN4BDvuKUZkrCgZNeow3iPr7jJ6q
vWV9ZYveydATFtT5wGqn1dA+i5Meu7pHBLIrAQ4FNqr6+5JqpD4tnGepXPwnla+r1RlM+pvVhPBY
PsR/GDKIC3NA84J52eKuJ/1X2W0dVRaLLqUHUGnNmx56fg1TIAA0ZcGD5U0VafVgiMVnr0BhffUq
sP3js+05knHAhHHfgYXkZQH5liS0MELaTpwMWXk7KhvUCcJqBMpYmPXNYg0QpMrs3+eiQvvqL/pV
J9r1ztyUaTdkiCETfB+8MHPa1A5kkNISSNuLysW+79YuU5/x1a9R68z5qTsuEHIEqz7W1XsJvLJR
87igqRLPNbfsNSDzPWWtbaz9JR1pmwG7kXvUfx9/F3xXkFQtu5ebOmG6Cr0Y8jICiCha3Z8NdQxj
YIKortO2esqm0fwDgKjFWA1w+0UCntQD9gd4QFNj5zfKXDGYwlTJ5pyg1XakVoxdoeud159nALp5
JG4ibPdDZUrKQ5KC+pdLWR0A0UCCmO1dgMHAXxl7uQDmWI5qS1lJhxeeJmremsj2FMLc+ThngjLN
44LxAh/JZCZn3q2Heo/UX0s6xjfz6OyB+iPvAyTxG+Z/l32ecoUNvLqYojScdC30U8MlIqMY5hfU
0+6UTjnUS7+bmckOk4ZqR++HkP8kBAmNrnSflOeEE75ZPryYQJiBiraicUxKr15jOVroiGpRvQfh
dd/F7CsXasYSk20zACXRcra55gbKpTwLX11snR8wEL+gejfnGeIgkBGh2Le63+ouZfeRIvFk+c29
WX81f+ki9K9ekP4r//rUjKzUDPD1p5gHnuA/c6WfMSd2w/K+tDu7ZlWy29ul8I+vCJgOF+VM1VbX
Yk8/Jn9OCZhniUqw8NGzCnz3HMo9odDh3mr9oWMdhW+t7QfErPt73u6Z791ttZkgtxby+wXWRbFP
WUtXRKrsn3rYJhW9rdnellxFKgHGDiX9NbmHtOP/UScHmmywmqLf3U6jSD3M5FrK5IGVh6MfNIe1
LHomniCcEDcHUbzv+ZEnQnbmxITp1r/9jRNTxLXHQqI8C9jq8P5mZvsjX+ptykA7GgYvHezidZlx
anNWhQaz6O6guqu0yMD14wWVlsPNEduHTlmC6fIj3fJ6oCDVfyanHRnyuc9rKcJR6iyr+GWs2sG8
krTp0l3nQzrkIJtxsvx4aU07uyT4y4VaFbKx28zevh9W5luAxAo+w6bUfZrZHE+wBo4j+/YLWTRs
mKveh3c2cjbX/fp7q8Vfljgsg0OEJHpKlWfE4tSr7F+HdGWKGG5pwMP5j8YVof8rA8+9aIoXdZzc
lV2wAVBBuFnk1CQs+/QmJ7d5fKfUY8ynESUGePe/Wo3AA8dr8O/di6M30j9E8gTsHuPGD3/O8W1h
24M2OgFLlV8dGJsrhSQEv5Qj4Jn8drne/jmSsLfzzMSfGZEQG3SLayubZ7z71Tm52CftMBLbJk38
K1/HBE3soWs/7aCviw4Vs+lSD2BwDt0pJ+cT2FkHH1GMe5bVzQcZDRrhWjozOaw+EKFYgtR+jp3u
9yIf2icyBZlbM/gG/IKpMMBz14Bw49B27sB6iqdOm7Juq9WElI7IHEiCToRdT5mjo2pToLuuSqFp
Br4kkhwRU6jK78T34BtwBtQeecGmtWdJ5F1TuOcv+Q2b7hXVXuS64AYlZDsNcPfVln5fz6HFTVBF
XBIULnv0KbnCLVf+82exv9N03pEK2JchDNFhx7SvHIvJ+LiaJyJFAxQwzAysasHj0sR1Mctqjaxv
n0M5VoP0LM0qsxsD01PMrT/7R8rdFC5SEe5xY4JmEa28q3Dk82yVfCyVMkTiIvFVj1pSP2nfHiCY
kleSBis7RUVtnGZAI2P/GTUj7MmryumUe/EkKUubugeYjXeKZOTNR0nhcaJWDSaTii8jngUYY0z8
x80soy1LykgJB/6DjEctB//hbH1CAhGObdsft//Lp2FTtDBO94BqcmoVV/1PE0nO4kK7IF7ve1/9
7AEZZr1yxgaA5kXq4sdPgA1ci7NhtKo4O7DAPS9smy62D3it+Qzjr4qH+RldOx3cvZEFfe0fiRxR
saiwe93Lvvqv54TP/0yDWWmeWiKyXFW1tCt9TQOtT80pYSjzKBCLvRMhxoBMj8/jRhoWvU4V0kGi
qiHAabcViG4qsE7PL5D2/uuK7CLhXddIQ7XsRrLOt9vE9vW/JyfGo5p0TkBjACJkGR7x2a4kwqBp
9J04+JhXpbBqct9l6U8eWnQaGnUche/6n3fz/IYRyMi/uSUgWd3TDwPf5rOu98cW6Zv27XHXz4Jg
m5Ot90qgqNJZLnoeQ9ka/SqDXHRQwZa1AkAqXsyfNXgQiTPZwMY5Cuv90Glb7ys86YrAJsrjs/3P
D+zjubxuIGt/MFHpE3z8Apj7VfVqelwRl4ULc+eKsm16OooPaRlj7XtmUKZkai/cQGdwmVK1reZO
32JmeexHiuydibGa5XY6T405wB1PiwxQLMf3k1iBysNeEpEVgOKOFp6JtyzNCtVcd4nnLxobHvkS
ZcQUy4LAFRH+vZWNeF0raZLeVk1a4yh7MffmuNzCSNxHrEMIkkNlUP5TWXb//PexjT8AtyZUJ13R
1p/2MU+pH6El3xiNtK/JAsScehZC0Uni/lsBk5AWSaMeoqSIZuduXmIl/kFau2E9LpamjeQ9NOZk
7oBG63EydcgIXx14ypWi4gNlpNq9fmfOGXx5Ui3H5ruzP0c3yxFgaZ5gnTNeLEiMW17vIncH8Iy+
6NT89Kvr09e89IwdvXIUKZ1ZUD1BVR9t2SYCkL8xjRWpU1qlBEjs9J9fKSdS9KZL+RVF4BX+I/LJ
0e7tNNGOfJe6Unc/Lk8JwrQMdNGHXcLe9dKz/GTJgr8+7zvjm2WJHrUhh1NbSU1KVzQGzsgwb58U
eUUzCndRSm91/bacT3g3tLfJrmQVDAfNRjDsfgLwL8hBeMrSWiCteY332TrBXiUO/4g0tjefMc7h
TBDzo1PSAGtTrbKgwTrXPBkcZEr3ubGGeAJ5JL9rpthNgYCFOkUBXN8UpvOeeDDnVkjmlH2NnZLD
e8XbSpWMD/HqdLli+iuEn6qX/wEO0MSvxp5FClXWnAgHwfVDy3ScExIDQ772J1Nj/4ehLfftfFvn
b9fpkGL+UdNpb+acRFc8BCqdVyT71F5L8g4qDiixi3UFg10GjoH9lcGHc5QWnURIgFLu637Mxe00
X7mQ0DE5IPSIAUChjlLX3t/BsgdlW9isTyRhz4gze/qKR72oZF0BAtmMJ+xF0ecZ/Yd9UjjZTuPO
QIKM5vUl+za8WMBAW713T/ELHfAmYSyEiv/rSGBJATuoq+fBC1tw/D3tiSEy7r35Ut1AOwTJD9C0
CJ+L4aCZID5CJa/8gnu6B5m3KiSPBSwDtzHw/gxoDBKg6FKDpZOMdTqa+JyrEE2pJiUDoYnLbxyW
ru9clqFJJV0OSwXa36kg/JvH+ba/yjUcB2ON6KtSCpn++ivbqY5XMfcTtK/WStH5aPhTiiR3bK6W
ynQFgFjGe45hiRGcjLcCTGJnP3TlMZZPuFdw/M8L4IgN4h3z5fyXq9Mdieh0QIR6JM8aMkb8WuhY
i0j9JbIupp3PeFAwV4kdtvbCR5oLTN0xyugwcr8ksU50oJloNoO1vy6SfnZ/ySFFHXRYCzT2ZbZ4
8Y31bO9Xg6hFr7SvG7kuBAcgzkgok0XpoHV3QQkJlq3kfyCu8+s87DRXb90S6kFN6iOVtBJZJgBI
zlZOKW1wMjxeFwGqFGXj0NCqceWjWJ1S8afMYAQa5xvGMlLINexYTlL8nEfY94KRuxLd6NaAWqCS
fU5gw9j8p+QT95L+lS1l2K9UUBat1qzvFC7nIJODlL9tONl0+CsT5+mFo10hmhm3g6SmG6UUvkZM
TGivr2Iuz39vXQlJw3cwBD30lREEvtWEPIrR0Vqjsg+5X6A4JwryQWyNqlprFrmJam+WUvHYx82N
MHxZx7KvYDjjm1JBrz8x4f5m6vFxsidUxxNbE99h7iZOJwgB4lS0bzcibCVGaTZKU34iqWtjTCIe
andzc5MW2i6fHom0LtV1Um4RLlVogMmcjuaVX3p5F40HiJe2HXop8kFW0peurWRZB4EdSm1pgvG9
X5sEEVXhE/75phuY1/6TkiygQpIloP+v7/UsM7aqvchYrhiUAawG6mJNxWP8e+gsgiOJZkNnAFis
Drgc4CuwawtVa5uYFOygsQpZlaWRbIW0ZPb3FzlE1ODY5Nk/jbS7T+DpQ8u2U+/y+7fxshOXyz5N
ewyhxsIuyQ+wGJlHWeLcjo1Eo4bezY4OHvEmhhkbx0hwAaePBZ0eavOWTrX/PW+xY+n01DP1hI6k
/tCL5v415wt7ox9wtkyqbr5BOUtVMuKkog0Y+KwwuKmgbPIxEdY8EtMIFVCX3HDCEMfcK221B5l6
13E+FWFUvqHSOzU4UH2+fC9GMkVYDL44k7o+V05FUch0vtVsJBbG11GUFOh1WJVFrJuE4kXoXTgG
YN5ogprprXfIJxdIw602C8gy0HdrY/3lhzhzEt0VdnSb8zetGEriltjzcB2k3GTJhKSRBbFcIdVM
8TR8LpNgd592osub/dVzFy3XBj7+IU/RfoXK3f6ZF0/Mh1zzEPnDuzFMKkdk1Cndq6BJW4vDQU/F
oRKwEBlC/MGuuwyUV1oRDeSpBQqsQapXS6FAmD8QrhA9lQi9B24BXy1WQXInXxkC3lDnSSYpUkuk
+a/G9GtXgyuEG4jGVwI9vOXvBZ2RWcEsrNIDzQDjQ0a7QVwLBwvf/+F4VSzUD2ywxvsvxWXyzlew
2RQG0DMfFbMkn3aUax++8mrGdrDXO08xZDDME9RlVAcMnMr2BAj13BfdiZsuf09NxaxSmh5Z4S6+
iZyA0w8VQ+4uEndBEn+awUFoRMbOMyJduySOJCFNCLlKT8qHijzG9BXLL7qQ8GqLD7HVB7tDtkxF
GLc+k6cvl5Y1khHZMo5FoKvH2fnK0Cq0NmUF4o9bvxd140KuHNWtlEZ1DIWlFZp+8IprbDYmOyPa
IJjKZWz5sXoWC7dwQN06eSEyA7v3J9VGpc9a5Curph/48D/3K1xZ5fU3EeDWS4ddHs5ST8F8suvc
2jVqfF8dPicnbnlGsShrm5iiKIZe2mVkuXxFmoW3MAGAl9Grw/05obXug0rVLMxEl3bsyZSMFoPu
hujZvD8RWsICMOKOqkMu4EAkJ8U044/MprroTBDNZqBvzvkD9b+TYZ4bA7trx3Ig4sxov3ktrcqN
+g61qB+ZHhseHnqF23Nj+MXalID2kYF55vHqiRCTH1uqu2in89kRG6pytOnDS0pmZ+S1R1wfmjt1
bvS7UwiE7eI4FgrFpmgi/yFuEmgUeDXA7/RUc3RqW05uO9pq3gQvrPBp9nao3inyxqvDYC2jM0aV
lQXeOUpLOd2Z0S0B5R3+0ds4xJYfZtzZQdCUQsx6Ui9wWRLUBHGOpk5G7kNi2VtJTHZiC6h6WFaJ
Ka7h1IQRKonERhmXk1EjhkLbAWnrCIsbbH9vCblyZAtjW6h7Mu1M6i8A1SqHEcAAm1Q/Z4aoO18t
KzMkJqLtBoTbZknkhNe5ptBFVFlCmxto9cXxR7CPHOqnWFCrTSPrOhtft4+v5eCbQWT6dLWOGriQ
Q32YDmKDM/wgEHEllpj1S1V0nhUlGbXqGxVWGe3tM8V8ysCls05D1a6JpQbsGD7DTkAjfm5qPcJj
ECQoL9RbddYNDOKoVhf6Usu4AuXllMBiyuRq86jZIy4EfY+DwSHEmXA5yKYDHyhYoh+nTeuxveLp
33qniLGk8eA5P25G7U1rFkpLxOoPSO0vZnf/YO3WeIiWV6KO26P1Nfsb3r2r5oK31uYGRUJT2XTR
r6T6bUof0BAVR8Qia5JHxJ+hbzjMMr9WIs+4DPrwQM54c095tFnrX+saqD8Q+V26FfcrbfhnZ5iL
2BWvAfeHM6PondujbckUSrLK9+cLYJPhisjffS8S30nUWuCMP6sBP0NBz2cheF/u0ANdcio8Janp
CrhAHj+HXKZO3S6Irl7XQEOBL+ODGGVfHqrA8dtlqRQ+QKFQ47HnGDioLcs0OPw9hhkNJcDUvIOn
aH6mizGCESqDZ2GnKeCJe5V81aH19DVd4lQgfjXCyUNcFXEp25g/lBYTf9UUEEWb1Y4IGQbpISpL
Gn+uIvMwp0W9uQDy63Y4zCSoPoylqtETgKg0XbNtvHNq2TTYYlM1ByGaPQMi1b8Be9t8VmpPwsrK
JGNiWP+LG0wRHXUTrMDh8CNUp4emrp3sQqXZRekGJCIjljgL73YU6J8OnUkHAN8p3Vqn62dZaRAM
lu5IznOeaDm8F9Y4wOVM32pUo4twRTPWIToZzprkFjebFvo47GrMI+pbfl6GBeE9+3YRua39zaJa
Vpp+t6lvutAl+sDqumdKWG4pqNoiKqF96A3kPHsr/at/gfjJuI3Lb913IGITwoRYEUBsY8ZksPZ2
3b4yk3jh7lUoDYNgbLSlY5CBMH8cVCfZYvHWFKO17MVSmzFuX7xFQH33qf7xu9+ljRC5xhjW6K0S
cptPkii0rsHeSpNHZETDy71tAvYY/6KjjoyI72fUazHvcQCJeNVdrzDU28Pu0ANkmcrjx05612Ym
BRWKPQUN/uTD/RY9AXaPttXgsMoKf0vfgIdITc2n9QyH68Bpran87oia3pW1sSHF/r04P6jIEOMk
S/Ge++sbpQRv+5N58Hl0Ef5ahG/z8nK3Y1PylfxZe9hF/l7v0kDrpl/iNwiqljiPc7ubjQzz0LlX
JBbZGDjWlWOZUclBaxzDAn7LYXEQHF+kRbkB+znUHqCDpI1h5InAFvLnM0CLpx3cKIl+N1UCTXKo
f8y2fYSCJTPRhwOoIIECaovbe2InUlE48+xCoQ2YhPZQxUqGy4hkfgL2JUHCLZou8EsuUrpQAVSj
JPaFZqWurNFPSoFS3UrBBpKZSY5nmytnz3URyppYl1yocGOLg2iIG73SqQBaubgVYfqdydQ31bd9
D5fa1mhvpcEzCFZ59x7+xsL8trYaUtZhso7IPYdwJoDYyRbKiJJRUTFKL+ptwPDjRq72UFy2gzgp
scULf6QOwC3CyTrEueuZdfel3gB6o74w/OiLS98mozkadLCM0OFMsshO+aSW94pk0poI40sAPYGo
pRJCH/F7vEctEDsznCt8Al3hslTIVkJtZp+FHdJegHOhcfxZ7x65KxTRU8uDpm5IiO5yNgyIEeNs
aWckc5RnOG1+ybHhaI+RiGwm7pRfqOkKHo7n003q2aBtIPcguEi7bg2Su2nNxWtlo1XJyrpNSPF1
Qx+yli1mTVaxOKIvaQtuNQ4VYxXcrUPbOkYVT9dHv8SKkU4zlP1Ul+ZkGxo/ChPrI5HTyj2qJzx4
wsIOD4T393wvzMqcKwIat2YRpGxYJHKVa5UpyM1yCH58fKbpfzZdhpzVd7z4FB96Ia9Kjqm3m4V9
ymYtCGbk5QbHDvNtWm7YA14aNv/DRSvpUcarovqT39bGQ0xJ8E6h4qwDAp2qpxI7vEyFRByYvMhj
sK2A5NJo6ardTfBvpnbm37L5W/QQlxN05eKTUkCmD/hJvmACmbcc7Vehc9QHktfxPbo+NhcjIwY+
ceGQAeOCdXsTUoPfKgUHftFux1StykFuXUIFuY7Fo2YJvl7E0POC/Z09ON5dD8Qa7pg4S+Ba1yvq
bPlBXXPtAYp5EQOp32ODV0rToMqFu26tIjach+jJclRkyC2twfSHYhr7G90Ronb3ARpNe+ykDOJd
V5fgFohUUoFYsZO5xGAeia0LSfmp1GGBn85hmkZtWuk80SvFJ0kuMvb7LnIH1FPvpwBQELnvzThB
nYAzx5Z+LWbNsGQR04zWl6fH5SbEdE6ZKGNtI9lGzZizinHflVU1QZ+mzUhvJsY7zW5PFBobr6qN
SCWn6R3zs7+PWJUrqKv6Dd24ZmwDMCC+wEp2JvSQ0kJY9EJZ6MYz+ZShPXbQLGetImtpRHo5qDPb
q6sqsR12i49N7c3kfMZfUNYWvCTX8JhnbHsIuBm63bcEAwjuAe289hhhXr8XqV1ECwvJfPCE31aZ
lG9pRiAYH/Vh1DexX70z6mI9p+ryIzn0qwaD8a4NHVTtWpFMtix7gou6DvstVtkAnWtHSljPGf9M
Uju+RMLq2ju7AhPSH2auIHw7BoJ4ESMEN3mA8jIQ2MnHLfkc+YrUQYcDOYS00Td7HB1gIjYV9RPa
Mfwk5VvmqwvNadqvlAFnlCk0msQRR27AZ7rC8Vi0XZg1Bn6IbQYnHMto+bdePxUYOpJFwtk/ac/D
PnKvRm+C5GaGS+oazuQt11Om5VRv7PxBKI9R0T7q4/Nqkzb1rMIOfX/sT87vz2KY0Mi3v/EAaZ/K
bCuP6ovgy55ro/gQ5/Kk4mqg8IWhgBPDvdVhXvRS72POyZXBFymeBdihCvcpRweoizl+ug2FWWZj
V86vDd480VZgUVKPpFYPyBRLqoA5PY+R2JNnHtNEJwLwELPuY8q9JYmiThRiDrFkFk637w4YNO5+
+RMAClRwVAHCwtsniBN0MAt7y7jrOJfgl2fZpfS90RrDBTyd/8LTD3bQslJ9jkMVq59rEw7S9HFV
d10gjiQAWwopVPio/e0EEKWAmLCGZC6V1j6IurrrvfRO5obwpq7gkLBvqHQPKn1jqkZalwfL2Znq
a0/0n1gKgG8ll+tmhYP34z4gx2EuPX3josbB1cSdMqRCtBHHHqROvy/G1A7iZlnRekyqcJAn63rT
MMbrK8FIZYxv8INuIrMDZ7EhVpJjV9Euakn9IbTZ2TmO0hAwa380vceczRoqDfL0xasKcFFA5rVS
iQdrWqeFbpSDGfftx2xq9ZXDoW6babdVsxJNp1x/SNDnMTPlW4x5gXOA3rwAITQVb1Di1AZEFDZg
IHCzUwwqW/+QvaeIMHK1/ZWZZBI2aTnOYTEz676MhdSBTfSFd75cUb/wPM3J6FANSkxC2mnC1cux
wKkfP4nvxzKF8G2dALErSHJLZRZWwaJx+ZW62IUQRRMETzUIHpKNoyGjZQKhJjKCyvegPVquSWks
my69abwKXRW60g93QFy5T/zBkt8MPu3yZ3V9NSAlPgfB1j39Uslw/Cjxh0jcLg8nIJs/jF3vedrO
K5MTAF6zzvot1U13uS5Lz+vC/VNxBeP9I7+e8NVVbFJot+HRJUMxQBJTcaoRE0cEoW8JCO9SZiYd
sbFjHWKptv0+llH30xodgvXyVIgErBer9S0HqC8bHlEZ4+nzBSLtJzKHzlkowoYXxoCd4PY3kdel
TP/5wvhGH/1HF1Rtvkn9L8pjkC7PljLmw03OjObaY+BUtuTBRWPPgxCDaH91avlM6G9Ntsqh7DCh
VKBqqhmwXJaqams8KdVPQYrcMdSoPdoHgROhGUYrHnzlECZHJOAax2+97Mppax6BYLTPGWJxvHof
dkrhnFXruH5vmF3gMCiMgdpuMY7ci9S3WxHYnKyinZNYt4jA6ZMy5mRnqO1Fq/gvVKQG/gyipNgv
NzvuQe/jD+kpkmeleJaQHMPRK8Ukq9OLnp244Se9D2EMDoNk2aRAslThfK7RvRNf5ZIlxbjP03qO
JersdUWbodMWfScypyPtBhbHH/UUJi1dEUREGLDPaV7C7NWhXYHsVgCW6sF93VZcfoDR4iIMSMe0
TtjF3Dpb2Uw122s/ALBSuFt91F9dlZfW7NOlztBSXh1EZja6hbN5vLxvOnKBOEIA91PKmztcQdNA
sR0aMC7xOzCzZsYhbYpPURN1dFQT6nEo1GiXfHdXDhGmR0F6sMyBwC2c+5/rUVr9rhs4sdZb+BBB
pFzEnekKk6OBSRbUr0D9ZaDRz8EIujz9GETU7fM6kvYU1SWomubgRRHcHL08Ayctk/GZ0xFfor5r
0XeaXJB+UuPDkSw7Q6TTItDQuIF6HBc9UI081iOLZ8OCIQWySMe1SCanpiWlSrv6YEoHEU9MBViI
QvvhYVl6AAneFHqzcCBRNvlJeDR9ZNyOKq4B9mGzYJa8+3quqeEIOet8N2JeIeI22Hujl75OT9n/
D1pB21jvkfRaCcybGwGdgNxm9P5+NYoHQEJ4+xb2GiUH8/0POV1Dp0SE5ctNEkqJAdbWJVgYwDl0
WhlyDzmonKJ9CU2XxKU4SXmxUb3yNXi3SJbcuXIp30WRTPHYdQz1nwffNBT1gA3pv0AI7MgnROui
gCUGAIoArAjOjHdqy2qgZBEwuENWKtwX7Gd6HkjkhpZXWQMckKlfOIigxsbTODX7weAHe0qGCiS1
N+FiVXyXd9KMQOrTKrgZ/uYO7LNhNSSQvxtD0Vc8V77/Eg0x0Nd+vcQzgcdky92ERYgUopwPLgvc
bxF2Itu9maE16xyyM+Xll88bjYOKH3MPKMU/3JenHCps9g7oRe6M4v6IHFPPzR2bAPIF4A3AquhP
a5yE3zgIcf6/EfZorCTcwNSwFmyZVd2rNrN9wx2hTUyy7V+BEfW3JLWp+c7ENaenoXl1rlU8Rc5x
tAYhryBkben2LAJu39waJzDNc8y/v9anHWAkqo2AZshy4thbt8XZ+BcZd1xcRoOFFADSuaGt3AWM
W2k7uWq9Qj52kcIslkNRUu+ibICYmn6SSvEfbTEahLTSdGPzdnCJk6Rm4a6MvFHcptNqDh3rq/5b
SNqK73to738/S8pvgErBn2OTAK3LiD7YWi48b7yRlw/q1O9k4J8j2ToAs9NQxm8huAzVmeJOo/W+
NE+NkCt0R4jAqE7SwjgIS6MpK4G9imfADXTF55cX+m84xt7Tl8RMJmSuS/83d/WiI3a9Rb+5N5WY
azIKrzIc23PKO1UB7kTle/AAu1ukFDGgPngChsIBqwuLUESjNePH0rvMjswNjuqmWRS+OcC3gFb0
q1IpLzQNlcs6vykqAUGxM9Tiu1PzV/Xi/T0QwZL5zb3vkwlBMT/iG2rulET9AJk4lLyXBLsr327h
ziw93YMG8NiPjeIguVp8V28ed8za7UcstUHO5EwyiPxXhVIoFwlu7k7qGMhLtcJMceTsXqXwSL1j
ErNniv5AhGSB2ouR0F/KrNSTqE16r6g7SVIp53fgZz4AsO9fnfsIpcr9XSUaIz7WOH/u4Ms9UCQ0
63fpZsm9Gqm8gdDBM8Iy+gATnC2SdEmdPvqAX9g+UvaKCyXTizdhJOHFZFlzCzOT3OsMZSsw58w5
QPeIsgnxq4u/qAHNB69ud8DE6T1MPtt/DS5qys9miZXa1JU6NSCc4rGJqqf22YrnGNRzJX+KrlkN
Wje+Wr36Rh+IZCuSUajCu4wYxQLySbB89V4y4NygkD8JO8l1VpuG5Ly8UzchGzgMUJz3qvAizDxS
cTf8efDx7AIqHftweEDchx1tuNO4lpB0xBfmG+C9qcIJoW5BF6Llx2pk6waacHalCcM1WZhJ2swY
6VjECBFI4iThK4rw2eXc5gV4TNZSbGqM8pOsj7WBACUMfkCrsJ8vN7irIDD7Z1fHlfx5EdwBTld1
Zefx337XnHcK4WJuwMWFpHPdYrkBzwasI1mp4YC+O6CQ7GpOeDWwxjBEQMw3yRbniK+tITBDuueS
CuRmK/iEYOlWS7fFiMIO0+Q+WOgi2/vTmq123u5ZADGbUoVHZ72XiOvW+mOV1se9QbAl3fA/uCFC
d6jMa7OT1e1MorEwRW9PSEgzt9fzJf3wa6jCGpPp6PzyNuIizK0J4DTsr9wK25ofP6YsppttfH5/
FoIFZZvznHM0jObB7qXfrq6s6tL1s66o4K9431EKJ0kcKYy0JLl/oh2IT4i0OVFN36rJ4t1axgTX
O3GCo3CTuGBcOPnB+KEVWy9V8wFytnagZd4yZQYKYL844FAobGgd6l5V6VwrZiCppYR/BZzuu/VM
E5M5eLY9ytDJJWlR1RlsjXq177q+uM6Ul3HKm4SuJd79z+Mi0jSAyQhvK58gkfBUK12UyqwKLhHc
w8ZzZ10QU6SoZl0p88kHRBr//5J8Wk87n/GClq3AxWLYmhZdwZGgtEn29mifm43M7/vSOVFjm/6q
fdvjhvPOhwgcr7V0xN2PNmIjY9tWYRP2EEYeNLFk2KRVP15WwVCsI68bzHsmjRexPT8ck2YOq/ci
RKi9wtxgX5jdmrRcchltmaqkD62RM+rsvLu0JybfsiG+VDCxLmXtpjacG7j4pS8PhcdHDgCxxI+K
MWMfwTNeWr162belz27P9K/pewuNjPJits89Xu8mBXOUEv87QZJciZ7xWDdV+OAY4B07gFTKYjmM
aYOoAqNPC0PJKHdT8vE9gsS5PF1Rfa7Dkp2KuASvIC1HDxjR1PdMJPNJIaNAWpbcGKEY8BScmIDk
Ur8T4t7xB/qnxE5U4yh+utJFe6OwS3y8qxoEWbY+EcO77DNM4cflkAiKP5JkPk5xaWeb4AmXXgRs
fj+gw3KXeGIM3yAMvy7CkCIkmKgF7Bni87CtHmed/82bKtpMv1qabwnkkGha983qL/7+JROVsk2/
VTZw9KNVVwDfR8PC34gJc0jDAqhwjtOuHTlQGI683kMtyU2IQ+SXjTuNiWKSmN9DWGaBAkF+EMVa
PmbWuJeELTZiAnnSR2snjcHeyUd2S8GUxctzkPezxqMIl7uTw8DmorxZKD28BVqGKJCzF7xTqaWf
41qSOzby7hxK8jT7FZ3v5LsojZluP6PoNES3ThwN07Gyb2lMIN9tAOlsLFw4kR6mURGlwfEoM2xY
P0bXuRuaJV6xFnQZm78lLwbSvGbbrQwhYyRLNq/4fshEHcX/E9Bshev7ng08EwoAAkZumvvCGr3L
y4LKVELvArAABHfLryavAvqTsm2mdFF6hWyL29YFOv3Qxl+EIBXSyL6Qz32Q99BfeawtFUdgiiQO
qtwzA0FLinyOpkshqH9OZvYDW89zm2dhTfBDLe9vOdQMy1zKLYEdyxtcxbmiR3N/Q2qIKwvaMgVs
W/kw7RB06Yr1YPh61ri1bcnSvJRO5/nkV3M/GgyjxEsJwgZ3tmPpmQwggcQNq5fuu85ici8laAq7
f/ORk1M6QZIGuqxR3mq215+/BlPr313cLO4ANcgQQV9tbryDv9Bs6YGV9SQ6ypN3ExBFRilVQX3H
RWfwLuRtP/H1U6C9oJxbg4uKAmE6bgrN4lUPgVD9cP7NsBmNy88EFOSy4JX/McTyDQXQ0SWS+9CO
fk2H6KeilWUUYRhTEOnNdfA4ctNIAx8sYvj74+R1RfsMVQHpDQk8igi1B9YK/t4HWJPPgzfobGR5
DfY2jA0DD2Bn5OTNDdK5wrs2eU+Z59H133ZGXC5N2tOVAXbD4+kCrfKpepNdNmXrGhLYwPdOaazO
sBlTbZPhVrVLH7VD0QIf5ob3VFdNy+32SDalbiFHvp0hiWixzYcfZWOfEElTjFzqpXT1la1RTW29
QaVzaRZglIkawx1Go386WxjwldyGbBcCC7BC4S/Pnq1eo96sQ/ucgOFK7cIIK17FR+cCbdYAjk7p
EweGWatQf1XYphnI5o6xwguVkuLVDP8kPY9FwszJvB92taomypRbb/OlQriXWLW2xxeAs6KLEmb4
Tc3SOMnNiOkHaoUPi4rMEvBmqsRSQbB97noPAVyN2d5s4OpnL7CLgpmAWoRlMowTsET4VADB/Hi2
kkbPqUfWs9js8J0zuBRr0eLGxqCH55zaN+8fTTO9IGZAvvpjWJVMm1zz3R0qa62Xm5z3Doj2/rbh
6yEOsCXkCGJsDra2VYSlqzM5ZPH/B3hTkapsi6nvhBM2U96MHB7Uu9OQqst12YI1sIJuvElfY6vp
O7jieMaR97LByTaWtXj+77N/tk1EHb8F0yJZIqWM8zYdv03wuHi5K0k5+r8Nw9fh4Q+kTF/oEhtJ
5fcb8d4m6X1KvJD92tqQK865ZE57E9rVoNuMC1XnWuvL952FYf8gvKIbLZhFtd1g7JEotIMoiYTG
nishk2T7dOyAaXLv5dBmZ5AOXqDCixsFrnJTHgUkq1xfkWjtWXt2DBZBjkqX4grcJxnltiYQMfke
txvy67cL/IXpsVyTgxI9iH9xzhrMS8G40QsIffa+crc+Dor0vmKYTpQ/4ZtUE3aa6ev+sA/PQIjq
8b653DEaXTtLR/IRKnfx83wmI2Ss+a2TsiMT7785IU6WhgmBkt1lsz2GeAdtPt80dac50qAv0fn/
C/DqRQpGIgcx73bS4mHrPXhjYT62k+tVhgRkVgYNHLl2hLn+GEY2/jN0JA5YCg4suwvuq5DpFWxU
o9egu5AC8hbO/32jrppl40w+4SvNa+qXEkeTHzG/PFfgzZ5uBwaY4mKdRIJXd0apyki3uZ4qYp0y
loAxWXFdm4Uz4FXO0UJpf5KgVRzPWpE1339Hzd6lxuIbyYlGK9bfwrxozqTZAgnKYvH9q48bZ9+0
EudvcvFii3sTMv3i05FP4tyLLhSj6CdrISfsW9MIm8g+NtiNNCOmTVMhKaC/9/Pagfqu7lXtnB0d
bDoxvNNtICTorlm57GduRRa+sZMA21CmW2tZbCdWKL7KBMXS6qxyx99YkjGAXD/+zzqhkWjIBblU
GuSlHaxnoeOhtOG1F4DTdB0UaKCk2o9BPXuTPIhA8gpsrpNY0d1EkmiNKe6u0ZIWJAFOyL72d5wy
X0mTypQ1NkJNXo7kEk1RdPvYv6fhBI/12tbb2t0BxhTKyiPRwGBbHoGxuL+/ZxRQQ84UEzGBV4rh
cvrvHHqqXVt39wdKJezBzVQ4IVNUU+y+h4hCYmEtJCNPyqfh0oV6h4LqowYmKNqYZciMJAnopx7T
8M9FFBG7HnklSD0LG0GN/p2466wHqn+sGmb3Dr3sqaWlDIgx2rEXUhenC+KIgQPRBr4NBzd9/vqs
fYNwpvvF6DhFo/DMmBBvDO+eWDd8J3p/8dxcc0bmyGE5SwftIdoKQx5Dhvv00WPA9HXu07lwR6nS
L+xeJ+G/FJRoGIVPBXblsYZ4YEvT7ejd9dOCILMa0UgNz0iSRRBJBzlRKM8S2jwygjPihEp2jBOW
TenDtjIHjsRnpBFPH5X9fYe1/C44QIE5qrPC86OlECR6SlqM0Qv5/bB//VtNtiN98MxMXLAAqBJQ
YKhlve72lVzrJVCxbL+Z2gJeVzrM475tkjudRPb272JEDxFK/D6BOIo+rJNxYiI4SZOYbbhm9H3t
2HrP2NQxkjdZ/tAquU6ZCrSy58AAp89UOTG7ijSR6yDwloPvyBSKaUES/VTlPCdWoffIRWN2OglA
7KB9vF7NlWRjXUEFM606ZfEINVQRCkSTyfhNSEEJWPEmDMfLh6gpzBGOI58vg0OYhDMwBrLtMkWU
bF3xOi+69UCsXPfb7rfH/RLurC3uN6ezu1EctQZL/18GR0anvNvBTkVqKDURWW9soNk0z4vTjn4Z
ZX+/Rfg+emgbai0z88tXKGHlLBqOGaOy9NB107xMhD3HHWa0UTNEjDzZNn+IDLy/UE304hL8rCmt
UJ8+8YpTY1b7LNH9Qd6AaSf5SK+K8nogjYtVVwVYxS7GQLizErSmHjyS1UR4wmFcEIWO7YPG2/QR
vxUMmgWTChbq+1JU99ebpUZ/a+TTW/ijBucMkvtGIqrEPtSHmWFjboXmxQuTli94nfVDZKjXh79b
bCv5NSXJl9JB9/h39tqFFRRCGxvhFwzK1LV6xNDnvHvAUrzer133X7g+/KVnGfUVngS1rDob4j0E
rSNj89dtpzBF09hzv2MVZsDbWLsc86FtPpqjOUYKi5Uq9a40UF7hSqs8kN5zibuX7LFIy+7gT+8/
aROzIJCLo5tz/d5XBqo5bHtKxAUdvo6l/uXZhKRSIPHSpvfJkcYewANyPoENecZ0r0ju7NAi7jl7
T/MNHmjKGnR0skOASo844lzrUbHG4IcBK6AiWWXmRV41BaOA3Sxg7707QrJIG0Phi9WClycDYwD/
VACL3KTNijGDvDtg+RNm2vmJsCbk30TaCoL6JXu2hyz1S/eCX35CUDFW75C5bgd2jjU0JrWWVwCg
DrvRElCKh2Xy/oVv3oOkvaME7HaTdsfrkOvH75wqQjeMf8ziHbociBaN7TtR28nLk5vRNrPC16PU
qdqEvi0+rqOG74/RMGVOxtE/aDzbmSfhmEezZDpPMWssjbuGLqh9C5oHLNv7WsIzdCpdkxGaY9FO
cfrdDbtpeTQz7nLlKZsc9geOoQzS7WNfdtq7rEEPfUNfK+sUUosayBKrfFdwQSlDx0aJRRbMWD0k
ORmwIslv8CrbHJpD3YVJMl9aEh0DggRZDOIE7Wye08AojA/HQ2OToDC96cTRTNMkQNfQ5w04Nn5W
efX910MPEYUCKwwhUHFxG8wZev9q5sMAB4L3CgJ8CQkYnSVHkx0TD5+/baM9oCEg6pur7y+W4DzB
ReAmwuMn2Dxbvznk0BQkPe2KpzFpK0ZiG0WTgjraHZltF28kGl38DTWZXvW39zqkQVUEn7V90JBu
HYGwvpbVX7IQVP0IlDPlj19dbi+IHfMM7/jhToaTCrimfPMgz6+5v2e6Q0DtvhZAuBtb9ZhHshzM
o7vKpbfHWzMz4MdrZ6il5/o5bTKlkHbhrxC+iUV/Ma+vQGmhgLTYjKUHFZCgrY8sPAwn+h0+IOFN
XBqgGNyPK4vIYM3gzuVCgIUFEmL4tSTlKQWxnyade+F4N+XGYnFUh498ll0sIr3DvLB8u2XBQiLH
PrEQJnSp8PXwpCNN3iEBtr3W+v1kYFld02zPj2u3kUxPjuA1zSLDDgfXVTEY1H+3gr5qbV/QJK4A
WZhZT3hjXzvsjzYn9FbYnDyttoZ3at0xDrsYsFk1bXQPGb0lnNFhJf/HRxn+AS8li3FVMtO6UeQ5
Eo7cfSeALinY9H8fCQnhVUmWhamXhvpnN231J7vALcF6uM4u4zUaK0xlKXxUcPDW/j6XARP2tT5z
Tt4W3lj4vRfAopU6jkFJ5Oy9R0mE3x0wyRAfKOeS0WkjKJYH79MLqCD0OECrvYvdkzYb1DAguVAw
4ITIkJV9Mo3hvMEoVD+QlTOwBq0somvczGJAie44v2b4Sbmf6UreUWdvAeJXch/m+UmVfV70XuLX
BKzjTU8+OBj4dQeD8Uu6yHjsoCcdMKJTM8AQ+CNMxR40ECkuDMn3pcRUT025sEdsgPxF/4jLIruM
gYck4YhP/SKNryhIRQmhvsSKmVSedLfRIvKe8nj5B2Qcrn+gIXMbnr1bHrxnJa1BCJqh1286QgrH
FUZPL3HOxhSM5p4BWMhA1xUIGuiRyUvkvb9SYfAGwLnBrHkB8mnn0yLM/8dxuSnuSFh+j+vywTeo
51uZzMbwUTev6T9fsnG+3VHsAmmTe524aa3dJCljaFJfbZxBmSME28x/a3RIXkEFyxH0ZeRu/mDq
uwJ+S/XCtuyrgAN4exCQpEy/eHC2iMNX8OoVIfJj9ajS9o3X/8HMxQPfNsji+QCP2cxibGzhNG6P
/UaG4mPd5kByKeZLrcbylLEVszCwxvPxzJ8qxqW7r6XoC5DhjgDiNOHf+fbSuxxHYlftrGVr8vNV
DNX+x7VoDMjQTqDE6NK3X0IdqCD1V2OiOFgKOYcUcKk1S8OE3/zJQw586Vzh4ItmrGY1IfxtWmwi
06u0ESHM47PzPa5MIw6wCW7d1ozK8jErO8My8OLTkOQAdtn2jgD3r92B2Arr9bPttywuymqkH7l4
kgRW0SLpbljLQb0Bhewf+JAMeKzRHC8rfQzRUNduCKfxkztyUUpPsMCjtAJM5IXHKQ1YJYq+flxN
fsAEkFc3X1/U9fLJj/W6xFZgi51SNz2BcJBg6jabOUQORWtzRogj5rG0nRZZ2E83Tvkrgpb/+/eB
c0dJHWLK7Xhtdmd/KLNxWyqYs1DWDunb3fDTEGOQLy6XKpwyXyi5HWFJv+25ucXjeajY4gjE5Gs/
gLSi+WjOo7s+G7Sw4smVuJ4yLX8jBkF4iwdQ2uHTQJFJfXmjCgJEJAhwnPbD0c4Djtpw/sju40IR
+5wXmeCncA9OMCoOux2V3/jBexAYVNHuc52BlhkBFnZ/52RzD/JtMgWDs59Ikw4cGPsdBYodUgpl
syuHuZiJh5RezNIeldJkOxtqnExno9wUpMT5xmZbl0IqU7rkpJXnbq3LQbCvhfdNXfmLo4U1KCuO
7UC7u0w8yZxxuXQv+synzJgklrpqhtCbO8buNzfWYt0rc+vjluTtMXoaOOXDjBjydAuhAP7Zm0gH
YUu07BOZH5XILed+gNG/nJZLRXcFT2XQod9Xp1MyhxIhdDDuHxYadX54r4qxSjBSvD+6DC/dk/Jk
VsLTKB391px1nD9pG4Lx6lBRVS1z1/o61akQkKLFODyHogG+JM8/hve16nQCjZBUyp4xYvua7AID
Ja3Tw/FZVrfhkGk7FN9dUlKI+s+p4driIBHO+hDYAwSYFr1EUL6WKI6q5C1ltXh3/ZHHZx5H4X0M
15oGQmHgrHskAqOnZUj7POUmwRlao1BBoP9Gifu9xP9R/TeUC6QB9lOdtU7DpoVvDBrfm77Y/p3H
ZnOPSF+IMATyS31fya6bY1SM36aD6YyVweza+xqEgj9knkQhrKgzIQSp1j0gGHLne2UJjVrs8vbu
YHRPOVjLEj21YV+zl+aHLni++UQjoI7vpKcx6z7tcB5850a03PTbujrVFZrp5umWtHYJcVG9DFrJ
4HHCnLsT0s2QBsXWyNuecuRKGyD1Bkze8OrbegSN1yirKLX8BdaMQwcxV6lXCdpM7sFcuZvB8O2P
5nX+zl2JKRmO2PMykBdUWT+9H+eAeyCz3jRAWzVoea8jfmC+/YpCsnjCLM0ZduNodmsoLys+lSPt
IvKCqYyvZQoZLCfvNcsDoIRAZLlKgP/FDvcZYpjgUX4Ejzn0RQsOm/38QCBZhP04MZEW9kPUx9hb
DHlUyo6Xn8LIc5CmDNZcyvI7Yi/N/hx3KHjCh5VbhHoMMCHAPW5hzPwx6jCTg7oqyiw8Ryo+zsvb
9lxMTfRceSM4Fc+ClT8qwdTUNYSyUONVtkQNS0GFg5iNKFqLcVQ3p8bm6Dil9If6GbJbSsM/dWVp
3cnjfa5W9Uv9vv7ZMnW+GtAlzQyb5j757mMJ6wcDdVbCCrvlZTbFaNBxImK+m5CUW2UDg2r8Y/9i
7Hue0eQMBfK+JwdzowY7qrLmwqlE8qCyfCN3SHnanKn0JIlfIpK6HTrhRaJ7FrLvZ7jCyQnNy5oK
nXQGCpZsWh+8eORcSKjjbl/aGAqbtQISnHkTRrmvWRAMVGpGRDl51FUIWinsViRpHoQ9l0UtDLkT
aeqBUZYgI0iFdMQfkJGyq6+GGFEydoUk427HffuPgvPCyerP7NOzT819NOJVlasiXJMI8QKzwLJZ
xMAxue+yKKScQuaZiJ/J6lb3b4j7r4Tj9NZJjLXANljw0wgrwYMVTyGnmLT1wxCSoI2jTRwYjB5Q
ERjBcBl2AJWeABawANa+7RH/8S1tpSHMmUDZ3lnEl4W/wxS1BdUPU54z+0osR6+D7EeSupkiPZc9
3bjhMfoQua5Pwqtj3ju3/N3P5SFsSKdjEOnHSktGyRUnJ16wcNeWDcKfXgkshNEuiAFRxmAtAXI3
2kqE/Ut10sGWLc7NFVy+BQhVH1+gVSCLWcFW9uNLTZXP2IVZ5hcBG2qkVuTpEAp1CMGcCj8A+UYI
wrMHZWLX7bSQa7SxE7U0gmjj0tmTIxwfdIS7Sqy9XnhtLQRCC+KVlLNTtXTy1MeT8dHU/d/I4Ude
+z8INpLQFgYCUgXdNiYuXw/s078DvdtQgmdYiWuS5OBLGrw/RqPtgIq24fQGfFr/fLhF+c9bdYZR
miq8XIz2/VhWRjl10XLmgRf9TtdMq833/Fox/PqyOcMCCoienjVCn8CAwp/rLwPU9Y0OpDTUsMPN
ZouaIvg8r6JGltzJsy9EiNBnyI6aP42RJP8Gie0F36/JHsd6zLNXF9+i44foNdccMziFYCRVLP5F
E8Y0Jv0XExNs/rq0g6gofUK1nmozOP2h4BKjR7nxqwHi3qFMJ3jhat6s/GCooDk5eZUc2lzEiuZk
y+b8fNI8wBUCB7De/7//Ktlm/4U/2x7be7QGtR9eyOu6KHvBInuYyPN2cmL1Kjlbzt41KrO3z6IQ
ZuNAqvN29JacND+LM4qDVPEm0leNjlgJSmQjSNXHuF+iznfn50dKJbVPstnxv0t5JjAgwit3dwwh
R9Uj9efqqWG+SFrfO9OLacFZIFN93xlxlOWRgYIM7g7nDBh2hx7vn87pFn85xOYp2KICsjNTww9s
PR/gJ8Le3bwa3lZfs2ExrcajgpuYPiZbAVvu7oTzhgc0Zlk5NFoPiNNNmNMg4bPXMfysxZosOV7y
YtV3MwEhr9nlxSl1lJhncMbV3qFAqPt/AXSB/nyyFwVBt+imr6pjUwkptJ1W1n1QfhY2pUf04AEk
bNwIctGUXZgZckY/391ycwnMbnF5JWWBhOrwqIOJy4/KRG5G6rZvACOAI1TMimoYhLheYb5EugCy
yK/gKgnZNgTJlgnsfM/3PMN5OYZWQpn/mGIfBWdcCpZV4Op5w/dKAgyfSzGyrUg6FxgMgAdBjM+D
Tux646HnxY8UgPhEZWFrU1+UNoaozmFSKNq55eE4nn5di5BJCfCIcdGCsKQLbSARO4q3zUfH/i/+
7FVVOYPNKNk+1HkcEo2Wo3yvfjefLx3tot+aWLYL2dir5ZjQNza6/HuvlBCbpvG0L2RSrsfx4ToO
GD3guxV+RWDKAMV/sVy6SRTrB16EJ2Z063S4/RST63CPI6uzTsfOlo9WOX9Nvz8zEOvwPutEFxHf
/2KXaR6ZXRVcdFUjWOgVMVw7Z+bkCFTjZQ4jStDwp5JeOVcfUArA86Q9ZcC79UqehN8UKRiMrd2V
eZL1/EreUbDgMNcRjwp4qTaH59aj5O6shoCiyO7D732dBXU/cnH67suDTsalA28v/MJqsz17Sw8o
muio1HR54N7nybDZrLtD+8E1C95GbKwBQge7C1C8GWN+OCENVA/N5iMnkeDy2FjkzY4BLDv4qhoZ
IQF9gCCZOuqjsWJ+sYwLWPwRSAw6iafWvaL6cvsiX5n/B97uX24kNFKdLf/AHWxkLGqKkd/AIjK4
c01vimP3zQPkXZX+sEl35TVB+PUrFGps7uC82b5q+l/jW9ZhKMmmguJGOarM/OFXn3vQmymijcjI
82NQ3hcDGLwPiVAFLYN9W/WzvnNq6L+2KVRmKLLZzS6Lhds5sx36G/FwbAGyHcVmutbFE+V+9qig
7eCq2nar+4V7HGF2vap4GJh0YAY7vXaclIMpnZuVQN/P1tmMNA+0If5wXW7QM/fHeBhE+9Uu7hkP
f5kdLfgU76keroEg0sodsfpPoBBqQ3p6bSjLWnaEYyXfWbYxqj5SGaKNW52Mjokxtf1ti+j4efz0
8Kn54r6R7Vl1F8JGkWRP3bFrgAu81MrSVDou7z1KNEzQiCOT7VNkACEy/PfSNJxTbNQ2Z8GfzrOs
LsneQNcwfLy7G/wBTXx6tjn6ON4Xkifv4CdJ3ARDR4ZS0Xcy4O76Af2fGWFDksMJdEUeLgUmaYaJ
EtJiCKFJh1Oxco1Vpkea+BXi9ay29leBgZp8WzsOye3kC4q+/I0TcGBM/QvMWEgLdeGW13LgKkoY
vV9EZtPLiaJUJ+VOlhRgh6qow98Fe8GcapiU7Lt7+fQHiQtSmBEqoexuvxoYeY6ftAprNFv865CB
9vXh5WUeXvRpo93DMChmdAAX9peq5FMnjQtbulzXg5aFaFL87cIcTuZU3HHAxZPqom7+IiNjE7kE
hTw9FSShPKWMhMLfxvEMsxRELRqunLCNv/3Ug2iwzdbj6PyCAGjVlvLedu2om4iYVnu1/QO4ByyU
M0GCkpbZia9leqA6uUWpFoz3VxWws7qdz5ztEV+d/wiYV7FExEk69TdSzl/G3FhQOmH5sHhnsqd+
EmjwKuXerHrLpQeXH9UHZ+9i1x0NkD0tHJSj2u7JsHvE13QA0YN94CYKDDubvn6hUi74qm7gyIbu
0STrSJtnjTGmE3WQ4y1Jm/khRc5BeV3pd9xpb19TvJB/w86Rfis9ygJLksuE+yKV3Bg/0bDQl8mU
UvEOcXkUJYk6yN7TxKNoF4HSzDPUzihAhS7F/1qp7o7ZV0nGkpCRoMrs5S6PbfWIKZ2cC/E+DTjm
4tpvo45Xla4k748k8Nt0T0iUzXxy2MdZNKi6uGFZCcqlh/bTPhnDKR+m+CiZrxMWnPqr30qG5My9
aUD0oWR1dfJ5ksUp5pYBxYolKGQ4PvsTxbA8Vi12H3gymQ9pm08sZHadmkMrf4TCYYukX8wBRI8x
G5USyIPl8pom6dfCvrC1PheBwlRddMnUOfIGQh/6Yirn7C+G+tv/RIL3YtBm8YCchT/p+mP5e7KH
dto1YE6uo8HgavMblu9Xor46OVtD9PG/RnrCQJagFpaWj2T4qOAX9mi4NFGRBYZwIfVrTXXTLf8I
uoPmTItF6J0z7wYMHsL+1d3+5tXKyeERhRIuWOgehCs3+HyjFdfPJ3TEvbT1y4TDAU/n+Y2JcopS
ZkZ8+UkdXTo0RYlPQteJDlM6XCzaHEyWMZhruoM7F8/PnoL8KPLpwKZVIKewidXlUZXJgSrl4+l0
/CR25RHnl6A3+5LtFkHSEyOjdj3ntTxPKxQIYYOjjmgDnMwsjS1n5UpiYl8K3lU9TfarOkM5HhN5
9iBBnyxwDiMtNu74svARvHs6QoC33pskusn6HpQul9sGy9ae0bLQnwmfJ5/kp7awla8KFyy5+8Jm
ReYvi0v50d0rNTz/abXWDziA/sIDGjcafrLnnm//qDK64T4SYOhbNfAVdrW5Md+N186d4TnRWzvW
gKMl/c3ZNsFsF400TQgIWOL+PQJd4d+QGKoaQAyngzohlO/ASeGOTKFgGCnu4L7fecidsZj0olQb
naeh+W6wKPr2H8TAdYMtoXr+YixMWbExC86rTqFbzVi3zmLQiOXwloFXWilk0WYjFxAtfcUCOVQL
+0N1Ra68LTY4GpG6pm7Yz7tMpKQSofJ8tFXxjdMwH73gmHc1DHG/prAg1CwiIsAANSQJeavLAkR4
LOLnXZD8EawbBz9VKorAcDEosnQ6y/QddT5cZoHcVJVOZ7i0ORyBTQQoysFieFf0xgLs2XNSADps
XELx6UOUVAS1Tdz7T4aSuA6gJwEkeU6zT036uOdjnARH7nScEyvoO2ELPCJVQdNcGkcg3q9dGFK2
qloyPB98rXritP2/Yw9n5II0QXZKVMiGBOVs494ICb9X/ty1nDPAkQBeO4LlgiezVUCsALz2zeuY
/BpF9/7ytEfk7N1gNkEH1cotZJSbs8YtcqRgOFNsK0KQg9xx8cd2FfNiovHLQaqnT5QqDlNd4QSX
nHCJTMG/gQE7O4M6JMdE4J7kg3Fui99bdXmD7+bCnQ8euRFUwPrSVWNvtx3USyYmiUTHd1McODlD
6wqbGf6N1reHTXXuSmm9J1utaQjyZjIwLWJznj+/2oupRNwVKd3FfnKlU39m4I4sLaBrd8QVxEGd
dNHSStM1BHmBhmwt9K2eINfTG1fVVMFJAUpNZRLnXWltqTDehbGXHjwqln3se0cBRZf1aeie0wzW
sjxX3AYl5aJX45UE7n84ynxiSlfNeK9pXKQer912ay82DHILI9Ig5R2UsyVAF0T8A1I6cz+vefMU
2zQeSrdB5NBGFRkT1GmUzUOVsY30gbTDDFxrngjesu9C1vihev+0LNQA9o4IjVcXU3Dl09oLaktk
wCP6qcqWKTpKZFyghcmYJUGgeHRxWmEVtl+ndUKUV9q93HZBmm3zyUajOMTf49lV9mxauZOEoqBI
yN4t1Q/pq4O3ODSnXukPt5dP559C3dXN72VMn+u//X4DiW7mSFhisjlZ2uNbjTcuitZpghYWNIkU
FsSzBy+7omOvQgzMy4kNW7or1pzUX+yRynomxS7ZYbsaZBJbT3XigONJyRFUyeDCrfgf+bK4VOxy
R7/kE2xHNM09FMKtpyjKCUzymSDRuWuXvsI4pHUqWCcI3ctxlNIw8IX0aP5GTRPq8JgOkZVY165c
WWhdlf6mimMC3qg+lo75nI8W2vPhN4AsEWU4xhom7b8UeBkAqEQMuFX9ykexvfoWalYxnw+LyDgn
bj6T/k1mBioKyMREgEc6rQxfJHkyaKVIZkd8D1+7AH7GvFRP4h4fTDr0g7Fnox8TqPMhfwWhZKkE
WfErF6GSjiGxEIZhmSjSZ+ZbjjwSp/dFTljiqwaz30fgWzQiSBA7cYkmN9LL4Lw8Q3LYtraxEiDg
TYP+4IvyKrpnZ+p7gMDOeGwcdbMJPyP0nXirQbrWRSAe8mYAy3n+TBLZPvoThpzIPsRYguZVs/qV
pyF1wBQa6FcxZ5+e72ryKg3MZTKzUBClvzL64O0fBwVFC0HRjUtIJBmPdgSzQxcTBrSXNa3SQ0NO
4ConxPQKvZSZzbgECL4uaUN0WMPGm5gLc5VuvqUVzTG98Ldbgq3Iew5ha0hdY2HgcbkKXrSZ+/LI
ZKD7UnUcGOZ0FydvcU2Z9EtFJYbRFK6pB2fxsDfVQOFMYnEUKGPx1sEiY38Vh9DbXznMkmu8+Nmw
nUfv9VhaXIY/QM/qaBtuRNRAGBT/wB0yrmKiYfMB8y6rWLvk7oXiawtcBLoBe6T7rfAf/ffqEslA
zyDdKgCGxO6XAKDodiS5giSWKKCy1zHH1bNeNz/gfriVmXBJRT5P1N50QBHSsFGm4FbWIFrjDp7d
mwvl7N1wv8T2g8aJw3ffC8aDops0cWNAPXmUewqPWJhhEUz393x7Rk2xcgjZbo03EDEN9cg/A14+
HthDxG7UohBA7Hdv4+Yul6LdfXIyxq23lE3tfrVTzogb54cWG3/Rpaovkf+nAC5T4grM6JuRr3z0
fn3YYSRIHd2uw+fqDeIhqFgnSNoFPg5mnmRQuZ71t3ZbftFq6uhZpBPPkf/EOMSHFZPx3hMkbCVr
ER7SOQvA5gvIW3r63OT58r2pPlSS0uLgnRt8fv2AvF2ufh3xcwOL2nAb5+IjqfDNhO4FKXYBXV4Y
VCsoADbj/VuxIJO/OMa+2skUHBsB2iPJthyIhcfKJkX3nha1x8dB8v7m6/I2cckYCdNx/Ml2DYDI
6UJapUs9Rh0hE+igA7J3Ty5p2K9mL0lSQRKjmZ+fJcW366kXmykB2I8hWZDEmH4ZQsZRFsYkVjPR
B2UUgSnw56D92nalcWxPKPFHxYvcd3p7OF5GJKhwnSDGR3Dy32MOob4V7pmVxuG+0jFP57RiG2Ng
ihDUdT10bdOKkAzdaFDqxRIqQswxxJZW91BwewMVwLRQlts9QyZ5BC0yj53GRl7lXFcyV+oQTub1
6D+Q7fEY/z8tMWuUONltUQx/f528cfn1Lwr0jwILiv1j4S+1BFAHBcDMhl94yWBUX5pSZ5ZhXemd
k5mGVDEUvzrF9fPFYrq1RRuqqtpxvj0522stPjmIki+6Cnri69u1sIX3ELTzolAR5g8EKtiIooiM
gC/heD8WKW13yguQ6APMCjMXHkbqO/4vdf9B5ByQeXdBnxJJrOGgI58bJ4W+6VwVVR9IeUSQ410d
QeWdqWYNOdE50pVw2pFYOl6ivxmJhbwrJ9EtROmXhvGLhhNn04pcaP6MBXkBHC9IypzTiOfJYKC1
QHmf0JuJvM3VbXrZ50QPkRDvzLQVRzu6glMUnuBWIv9cUszisummrdmpwk04SN8D1apkmFVrul/l
5nGeStDEMeVioIYN9Lgu/LfUmzqiaoJLR+fE6o3Ko7MmY67sUTkn7FdASodO18s7Zcj5UFB0WL48
icOWqC8UODxdwRc2eL5jJcHavswKlmlfaAMSIURu9bZlHiGm/Zifeq4sBjHh0mcaNHdDMKMq8XJJ
mfhownoVC5T6puNXmrTmWJZKyPKwKJGLy1W8COp+lMp6VqLGD+xRqkyyOvOu+U9N07GqjrBSFHFe
I+8pigdOFGvN+LJGSfJo5qiUqdIRTSBvVOf7wOc/EvmhdTcrfWmexWYVyttwmAjjuM4xhyxNeVhT
g5npCyhMN08l3OXTAb8FzT8ZLc1FbxOz/T2Fqe6lgm0z7J8ZYAP1JOVO0/gUnOFpDRNJXBmX7Ht/
yIjnG3f+QezS054xyecbWhQfx9HxxQtoLcVHa+rgtUzFIKoOHm/D2ypLlh0oG1sLuL4xvFUrPYna
7nqTiqD9XB1FPmSsu52IpbnqLNcfLgMa1W5pEPDnfmJUjLqVEUO3r+qRzNcXp/cVkHtb7MYb7jmB
2KCrlwIqOHigUVVwQsbKGne2PdAaVN/kY+skf5hFQBCXyMF7hIGvjKEjmcxlvKoAB4kdeXke0SQc
Fsnj0I1Lo0IZn6SNY2ro9ArshOKn7H9YGad5hK/+Zi/oIVVtjDfiy3DxCCXwQmK5E6ryx8Ji7q7B
iPHb1O22HbOQYD5/pAsoWTzUUTkz+5ZKoHR+9ZQ9JkFLyLvBqxWiTopjJt3PgH44n8nQIFPObgnm
5wTPvrGDpIx1uEFPmQVWin4Mc+wm1rrI8O5Yy0fgC4+/Fj5VByBG2QT6Eet5DhYj6UdeY3Z7nn/6
PIm6VfrtDxKdp4HoHzcT9LTbSrylfZ4YdX7o+rS4ZP59QzdnMFmRL0e5yVF4ir4dwyH6gwXjJgOZ
wiH7Wehk3GDSTHxIU9TzUdKDx+EAZP2ZqihGboVREG1HDaCAq7Op6ITXbtRdE3Us9jEcUSniu8Aq
dq1NUWi2blZBVWeUz2hC14r7cO453zA/32H+B+2wpLAk4kWkj1x+T7aj3VxnG97SGh6eVKEVAR5A
nj8NMA/XoA8N5NZx86/D/rGXHaMiN8rUQ5jDEyDfMipf751tW45D0wotCfHsmw1x4XW9yZ9OK2fx
KcDibd1HUZ+Ei+WW4XwvUXrALIHZsHPe6utOgSUAD+UuPfZaTWFdIfLPo4Qm64LByAOmIe0zHPzG
vB30pQM9PloFoGHFY54MolpRTvbb6ZhzqJAW0DlfoykfRQaLNkUNzP/D/noXJE9f73nOppEIzm/J
STZD0MWSexLM6MqJpcvQ1yh+BEUlRHbqq8FaguSFVFrfv3eljehoe+whkF5e0lnwwA62KzH7J/pj
VQdRXwNgQ84JXFuLuszywM1Rc+J1zp73lxfEyRRgHdN3XeJdmD6U/30LOGj2T30/BhO4hGp4iwa4
AC8/O480nQhdkkTm8aRpkCkNQWeXj+5VzI1cYUHLmzUa5ESCGudGQ6YsXyfCoANJE+E7xiH2a+UP
vZYKuPQz1qlaFRbZ/AMaqC3WL5+8amvtoZY5tUIqwTSgourMGvpwWF2CnO5YrUxvibOFDfhHQprX
YkZlRizjN0FR5eJFVr21XtZx6qBjoH4jZZfeT5eM0XacyjYcf70yMFr6aSGDCJaNYorR3OIVvVsC
93mlXxYkjauTyTNBsYshlF9xKPuojoRLyYvRYaNfWzsBz/nYWq1LYVx6PX38G1vq2di0SVsxiGg9
QI+XsdhCxXvcQb015CQpIxuOaBACZGoMZJA+ZYk0tevdW4sa1lsyuHvOd572o2dQa1CNEKBA7sWe
n7u1/s0HtCZwwyPgHElaz1bB2wh0/9H29d9tvlxwy8EcZlsllwlm579O7CESU8MxrGWE4+z7raT7
DYKvuNsL2v9DnsDGo87YZAHqkG3T2sueg+STzfhvB2pDzkUwRbPCXwj0L0J69CzNNzfg79BiFE7e
xg3IiJvuDz81g9DvyuGN6382V1qiRq1OeJsRWrAH1qdQjGfG0UWNMTbISW5OsZ/wFvdd9/rNnY+W
pyl8Z9lfMCAh3Z+rVuhWSw6piv7ZfS1CBt4PZfh3bbh8Zbg/Y5StsS0l3AT/W/wiAiZEsVmWgTaf
MDVtgCenlYSaEepzOot9xH5jKMhtL81lL/ovPFXeBhZSrlTwbJ3iIlazeAzIVTJtux1pzJH2Gc53
Vd7xm+KoUrc/SUNdEYoKPurE/BQ8RxnkIFnCFed7pJJshNdZeHPGHwzU+mq/WX8Zphdlo4QCL8ad
ijpNEbPNoJ+RNf/gXceTD4qYlhEUVsQhTBDFnvat4snT62bx/Tq04N303Eoz9CzU1b4mBL5f1O7y
2wqndSG3gd0bbz3sjA4S89GGWBD5OGKZWLvp/cPtAQIhyaf1z+uDkWI6E02zXwGW7BZhuquhlyxG
qEp+F4IeR29/TrldThVUaQy9RlVtNn12WvdRni7y53AM3QMlRtOSfnFFs6Qe3uwOaYmt3QOLjLFJ
S19WKeDn5QbJwNI9drll9Z5KzzAj6hXw9h4PKwW6jHGVJ7N4k2mvipyREP1wsm0rEr5wC8sDkUKb
A8VFcN2D0bYl+Pnu7NCjQCbm6TOuMdMgAB9X6zqo6KElvC9caI3j/ySTQGb2Y+YzedL0bssgJNg2
Cj/qd7tJQ3AttWDGj/pAvbhrFlR0vo6Ws8bEH0qayiP/BlIZ29t8SiRK7/UVkJbDaTeS6dhrno0D
YnveZnEkDeArP+kDjexAW9Gm7WdN4eMFcP2Uy1wpvtypaOVIqkWg/ArsDDLXIabqJTDUJ/EAFJqk
IJ0V/Wx4CU4I0l7XtCYHPgiCZH1LFUJIraH9pVN8hvGv52W/mu05k20eSrTKHKqLT0vGftkm+dWU
ImXSZ4Nwwhd5bQ4rFCFSXKNjFfPP4xWVsrskrGH3iOcGG48hZPPU9zLK0kCD9QGTqiyjZt0DQ/mg
2eVze74pUm081YyyhltA/sGuBN6XLmsBxsCFM+eD/HzH2K572CO1tDta2BEwosNZEmeEn6gHxwlI
ohdgpFi/H5YZfCOaAyUH7CCksIj+fd0AwiSQzWbkyeirpzWD4jI6nnW4JoBeci3GpIcT/CfEAVmd
YTxLDjsC5QDaWxACm31CZgowErgrd0/1EXFTlSg6IE6ZoCl7wi+UJeP0dGzBbtwBB621f97BrPfS
TXzfJK2KU+txS4sbfx8MUprIJladulXG0Pwc5v5W8yePfrk8JTFIi7aWvwGP1hOTkKgQryQVPJpI
UhRBnlKO+RXIIxvq6mwK9jj2t7K4dNG1JPtvL4LsrX+JX9FWR/WtwbawIL+2eOHVTrU6BtdS7Gi1
VSBXv/iQovu08CBZuPsN9kcAtiY8tvpBE4r9dIeLmssAtdFYzK/Zr2QIee30u7bZO3F2TZj+Q31C
4wGAJXm4ccY5gRnljHGbSuYgazlA+8MRYg5N54dDJV4Ch7t0RM3bqknfZni2BrVQp3oDD1IUY8/3
22CiR9bhq/K05ZRiaXNc1Ha8wSk82UPa9cjvx1MPKoTDhbKrP/stjpDE7kuI/JZf6YRZ2h2qdVTu
lmgZna8W7/xoLX/SdjQ+JLkiHKo7QQTYCiKdUFBXmHZNdO2RvyQKZnUVxsgfzCRJTPzcR0tSMi3y
pYkZ53+g/33bHxEvhAsQbbtQoushq/RGHJekAj6zl6l2J/DAA0IjAbPBfqs1hIYZLb+/NzGnezWX
Yp+N7N2Dqy/0r00L3pAa8REItjR1oeWU40dqt1/XQnErtpvhql3UbY9Uw3EO/y338zEH7Vj+l0B1
1ETugZJ0TPmBYZrStne1JmxCy+q/yQtEdCQOdKABCj8iAgfOiulp6//IizdKWYkJ6pAQVaoUEEFD
Aw2B0R6WPgxzmNmgpxLh1/IjXbj7TMCqs+grMi/MMaaLqP2bxjx+943ACmwSPE1RQ9invvhoN6Pk
X1UpJ5VzAvgIUwdj/UNH11ncl7CGU3LZeoAyoJeKix5bPxHT/xmZtrOV764ARZTEHFVTHQ8Q5Wyu
MJfDrTUOIzJuNIde0TiCP1vf5+jbIXgAy9Pp5STjJKi/af6+64e+QtbyZGyoLBGy8XWFiBR+ZP8S
gGSERjphBSfuPfSY5y11ymwrAEaXtYvMWE0zOvsUkrWBgwFxKYn3t1pLZl9guvxeVvbtgho3fRDS
K2NVhtetxIR07e+sTP0EWdLrxjPmDdiSu1Ifage9uvwfSw9xQj4FS38sZCEamY1U0DPbpIDpo6+4
IoRuKVkSoZssudGK8ZMwsvgB1H0BF8cmw1dH2+px1d7qMF4YQwCsX0Bept68dmyXHafdIOREExTa
Lj0LRGFpIlrEt+/66tjr7YnVEId/YkXeBJ5dqezBnNS78qbz67kneYe6icJpMXMGwcYVwqGmyDBY
ZUCN35ZCVxdz1LtmQ9ke89ieECs4ku3Gd4J3QCM3Abmyy/dy21hgwwlfwn0yiyomiRXeUOHePLM/
jd7rKHmboLK/ezmhAbHr+R3C5vkkEwIUlXR2SXJQR7KuI3mWIMezuW16Ut/6sKa8u/+tNEguAFbd
5TrNJhGDap+BhJcTCW+z8TefZqApXClCU5EI4yk8dOVED+RInZ09Nvog4rGweo2MFFRlhpNpjaD+
qup3T1E1a+6tTRVSuJmYCfFS9qAOuIRJOPKYt8qaaq8sgru9xJJfuLWPiXNyK+7JFeM+WAXxQe4n
FBg4WX3LWt7o994RDPTeNRpxkg763HvYxIpKB7jl8nfr91IwYKYYgmy5NFGMKvAxTGHgx3DqLclU
Bko4MgJCtSy1DXicdf3THzCykifblAEW1/dN3nMRk4fTMZ+Eq+sLwaPdYU6MqXtqP8Zyndxv4fht
iiq/rVtMA7HF5YjhjM0G8xXGVW1mt3KTdDmIwyCW3fHB15adOf6QP7HCxDmhXbVTdbMBhNqNIGKD
tEci16MfEKp9mm2AeL3jT5/0iGd0lBOtPMjDJyz8Lgxn7/CjdBUeSNQI3Q1jdXExYIH3TqAkHDZI
ediUcDVmrI/P96ZtqNK1bgdmjbut+3o75281Z5/pc8QqGNnFpW7OnFRCXb9YUzLLD21aisJgT249
ok1HAQc0DVLEFgJQFz2lVTpjO/OAXqOX6HT2J0DsXc/60LzdFLO9EU4txxBbG55Hxud0LMUiiI6E
sv3vLXAjK3FWFV4gzE4+KzsU72A2o18vfsMMdenTpFZ73zHW+WyaIf5lBH4xdUe8vJEOlUCtAEHC
YyhO6uq7cHXuVfRvTv2Oy1Apqd8uql6eICslUgrhtVw9nnGvTFZ/6Fnucb5qrU0rqGZ0fnWmHGo5
60pmLoD4hbGmL5JBtQDI+1MvpnmvHP1MvcuSx21qd68f8a583JnYksE7Pnf1qitYFxOR/elVwJlL
jHI5Veftxjj8rfb7FwJ4iH2xXvyjV7JsUlyCYwIm2XCOBnaSJwBR81txk1iTcxZcMBJJ2ydCZ+SW
yVGfiCZz5mRa85XsmnQceiMPVltvXttCITrTitdPvyM1QfX03RPTOMXSy1Da3wD8x3iCH3clXDGV
cIuzanIWvoB3qKP9P9NZrW3vK+2xUWPqGwM1yrgLRvNFO1B+UivGMxBsIALA/sgJSKbc8RX3OAxb
oV5wOepBbflf8Wu6HtSeV46/WHQKY4l7+8Xj/mvtw3Fi97GWpaq9zfZrrLd71/j5NdhG1U+26+bc
MN8s5lral3bbQttnSJ1qg6qLIHn5x7UCrs2ppxSkSOgWaIGEw0UAE3gJ7qhQO0BDRBpZ4NBVm3Nv
69mo93ksaL3B/fRn9UoIEDkO6RfajZZeo3PlsrhzH9AbT3qrFyoSHn6UUlNMp2rz8lW6/u/wd6X2
37gCoVc0RltYb+waz4ntNGejSwCI+hzh+CnrMEGGnR//22nwt0H9vAt5hh9DEgWJp8ZU6HTE3l7a
Fks1z8awfBWZQrhEwBYq9dFGOYyRH7G+jKSX3zGTSXckL036CuAKs5g3HbIp5MJshT8gkUF4YMRX
eFZwj0eidoqNkfKqRjUx9RM8P5XVOtmZp3aIW8tmCoQiTvol64oMUNtePZOaQ1nbGeMBjXr/y6am
n3dCczgMmzEyRt5/sN93gilS4X+hUZ6rhvoUHTuwYUipwb5BVJ4DQjHpKpiZFNDltwYDPYL+ZNjV
nGulj1fWNP/FYH5V9YotwSEzaEbl7WwQ4rXsZwCF2os3836ejt3KPdHmZ2IlNVDc7ihwXa63vEWt
5tDgOJFG2D9JkIzLssuusCkqAslh0B/e+HS0gWpheFZYBqItvcM1YdMfqk36ny4/bekecsN1QVDz
JHBbNX/AYvG4mhTMAwggCQk9XypaR+G6VR4sRbuze49zDECheuL6YdQzDokQ+eu6EQQPNOVnzsJe
TxBZTW04agSVHIzm/YQoQBoZ78gslMOKEYB9k1UxWArQxhaJEwDzys/AI+Q5jt0RW49kJD7vYuqo
zgvBtqRFF5KIqn6Lz4NTG1265LI7YKqcnTjeHDyGqE3w94loa+KlnvF/lAkUw+GjQ3zAWfizu2rs
5VQ2Wg+RvpVZaqtV4su8dHvW+jmSt8Pb1+aluz95Smj6fqMLjzCsTqS379c6XUQmje3tfp84Wcc5
1e4z0phEob4wkTEqKPzn+KFvNtasY0YPvZxXwD/OjYb8CDmV3bmIxjSshvIQFFcOj6s2VkFHNYs6
4b5KUrUTHUYT3h01uLVTNfUFv3u4NT0PwUOQIdeEA1UxKidDEp7VWnz1IHIqZYkwtTJRntRM1a90
+RByNX+hTlKGR2lL0bBhhoMpcT01DsmGQxdXHr7zSgEmHhujogGFGPDQTC/TmQfdmnAmCh0q+vZZ
RD3Hj1rc5InJ0phH1NmX7SOy/0DFlKHWv1AO4T5jQPClwQ7my/UyyG7dV6UeF4K3pU0MtQteZ3Yk
n8YqSp9Nrv42yCwg0Bc7GOybLGC/IXzs0QPDAFYbNlRg+An+fsRrSC7DI++dntrbVy14GLv/KqVq
gw24GJWrkfx/FjYeeQH2nf7McdSUEx0Xo2L6oF9Iq8c0XqDonejLvnViSV28D0x/k3oS3if5Ljjq
/T6saDZehjGz5VGr6WBxeBIcSIAPydwNvoPOlWpeYmeAOGStha4q3IM2WwCiLurvgCG1+nPvsLyC
JA8AMJOqaFYNF6ODmLrHu7/8RSt7gVh0mt8IWKYXAGAausTPesR0L30FWYdHqW4aI2fenm5uVEuX
KfnTLuirvjBpp8DLc6F0LzO751+Dp3zmeIkOjHXTcb1uMbtLhtoYjULaKhAwWPuBsI4TXdkZnEyN
yqQkSbzmpVxdDUr97A0LxTIek0b3+294l7h/vdj5r/PPtLYk2brWOFwgFahPNwuutTuinxCeUcvF
LFkPZRPP6dkA4wq0p62yrMizI7mfoXeOtMudUMhmoFiffyN1LSM/RApPtAhBuTKcqrkS4M63YmSF
3NIH0UFOGeP35DEfAt+ZR0btkO+iJ8pIbve67PBLT7IrVpIeV+zo60VHRqYH+c4Y0uAqv/6Nzmeq
vpgUKUAOIvWqDLjNw6Ksm/JNHan8UD3rc6y66DtQChMl6C2fVTrdKtyAN9FHP9HSqZLBwij+OHaD
4BA6GGzAl1t7KPFVgZEilXq17IIZ+/pzzgq3b+KMl30d9P0RGFLwimcQ8HPxfl/rciucANxaxtDo
p9iOTpufOmkaAdzz+UJ2r5qIpQdGP8x4iQ+ZX+0fipKsxOT0qRQRznjbM8g3TaA9OCD38PXxPbi/
N8oGbBLSvybfFu/N0gGWBuNFxYAY7YjJPOt03TCS9v00ZMI2sdhzwUvL5IQdJ+uhJtHO3wTh9a2u
MID+67lmkQiDLLeFcuQTM1acBCqcfSiLmcvZ1Ss5Hzerk7wOhfFszeBIMHze5wrMXWL/uGUIvvtl
zt7VzHMUSxRZ12yDrS4DT6MWWPrZX6o4EVMA/blrrIk49XgvAcAhZYqm2Qln13kDkfohbXNcl8pb
ac+g8bcF8inDTYlE8/oyP8mSuwZxcWp9xGf6Xhsta/F5CDCARz8qI4xwjnG8UNTXDwKYui+riZ6M
s4jTSsBnnvvhtMUTjUmsS2ZrXBpX6XSGRuCju45cT6y/xcSnByf/IX8NdVlpRsrV6NRCehi6Qei2
bf/M8BHq3/c3hOBBzu//tyRwzG/hC8wAjw5nFbwG5LPm+gHLJRyhKVHsK/SbyVKYLTh90qdMwUEV
sAHgfPpo/di2JShcFTXRM1zxYTkUc0QvIAaCYg3hJzLz23024qT3Y/4mXianIa7vrLmIyjSJK0mP
MVUq6cAAbf4xqqZTpUc25tsn4/JiYntl/8hmgaTnuHJuygah6G43kX20uFxlmtGy8doRjG6oCprO
WZ7OQYCDK2G41Hys8lOEIrQ4nqdqnXMUIzkGwC0DYcbJ1qlkds6Lf0S1GWpyZBMUDpJoBke1BEgm
/Q3Ljz7zYVkaY/tZKCjmwI7an6zv4B/c2W5SV8o4M18tLrdkZZ+FiAkiQlj+upeZlN2zy+IfncH5
27k6UITpJKPxvCsKPot+d/4l+3mV7xQ4vQSrEGOymCwubrGYpbz0NSaiQsE2R4vQY/lNjU7xyX1w
LfSDFa0F7KL2br7dKVn6zgOVmedMNi5PZhGdk/jZWTYcYRUhSGa0idu0O4vIvSb0zE7Spa7efVDB
rjYX8wPsF4YvbXbFHHY0ehYL4sNstGcb+FJIqOqK+t/Y1ixNY0Mbhmlg5KVFyZj7h8FQoUShoMFq
pbs2MozdyJ+kBMJVa7Hug/rOpwc34c6ZJyrwwRnYAksGfI4YpMtxkLgN85ftiVpEqzDbnPQH0FkF
LbpqKelnVrKd5N2lEvuyPI2Z10HcEZLsBgpkaHp0emsl+W7m5nCWnwaDWUFI8pAp4XEAoszKImCG
qZpW1ddv/v5cimqGZ24BBU/ou4Q8cG6bkquMEwBEPosMj1OFslnipPyvcI+S0d9eaOi6UiUCE+kF
20y9WlgKyvCek/O37+WsHe+Zt0viktxLnLkR1VZAaaP6HoD/nWvWxPAdU5tQmIMaTWeibW4AXLo1
hW5Rg+fWWF0deb1jK8zgKyPQ7TIL+QRmO0LNG3gzle4wWCHNSR5dmEP3CtIgSTV4vYJqR6gImxop
LkMGf4383aY4FMO/+q/3b7cKCyRQESgu8EtZzGWRtTU0SLhAE6mYbOfE7Uym/sb8XU9Z/t7A9L29
FJ1bBx9g6zOAlJ0yy11LfCsYrxkv29217ryMitKpsukD67ebJ0O4qP6Mrh5usRV0niysm7lAa0UN
VZW1Ia7DzvnhucK0rjW2K0jN7O7/cI+WSlikmN/QzQp3ztfshq2KicyXQdeFj51pvkAuclJoBkQN
8KKC7/n1hJGfUAwUhIvXuY2dwwLwIe2di5u6y5/Hahj5slFVS6AM4nU1VlZ21WFAzyKtfna/pvQ4
dyv2lLIp38RJL4Rd1pgIWB5nZY4QIbnTvizpScH2qukGTatvQ8+UIbx1FinLsbXaIRKwHSA74gAg
XYTMIf6mwT9Zns8v+EwIaaqCK9w3WwAXwNad3KgXUoYkv8zFmQXpenFMrXgk9lMie0eVmxm92xn6
RgFKZ3SUrJ3nh/jKM2PVwgU38uTeOcVm2xuSzvc6Nz2wrCbbV5ElwNmK7RBOtFlxMJG9Y68Y5N5u
oaIz+i4q/vfxZQ1EdCoztT40bukdELCcvK551G8Hxv3YjJd480jeZOIcmAfNEKVeZFFtKQhuSXxG
pXU8EQVElWGgw1UtoRNKjZJjhYEuP5T6WUW+eyO0H98Fp1Il4dRcmPmNSIo5ZNVfujhQg7XVaPK3
UlIvCa7sgd1S6D0iN+ag13iaTk0DIVYLSlAoi8ZAdhI+VtNZP0i9cJkDYqnCCQtU8/41wNZRap2U
wdzHrcRclloN2yJCw7FeF1G8hUDCK0w9zSGG3t9jTXCqhEbwjmyxbxuL0qViU0IWch3IESN0yCrG
4aQsYHIW9J8FDDlrLky483QqkUbqYX4Aa6I3xVlwZbFfvNln/1ZN8bJb6fN9iiE2UixijJMX5SQi
5xOIrdS7FNFt6AzsmJbiw6x2DMHWJC82CgV2MPQEhkR58J5WrAsF6fG5xDMSIl2OShbev4FD7Dpu
sz0vq+gR+k/6WUgU8fkZEQ7XZFZohlkgccS/L7DimoaEWzXReLKip8gh4uZgLRlZMB7wi1Gvg84B
iWHTjNr1HjEZzMoAsWsP0dEWPVG95MLmQVBFCOol5jBZStwK7l626jCbbU3UXUAf+2kn22fo6Y/k
ZqpjdhlWRDq7oUEDwMQNG7u+KP3HdMfyD04AZgC8PjD9ms2dYxkW+rBeIcHfjriqrZJ4oeEgGgjd
09ivLz5iQNmrZz6d5Tva0qaUeEkKvtJ2SKqr/INh/lXMxCbuzXWJ+Y/AhhkxJY5tOvl1xOXnMj9/
bB/AsgHF+zgLP8Hl0UBpc8vOikgof+PJNSYwpU4GVYORc35mZ3DA12ASbLm6aB8R/8sAszRZ5Wy1
5tg8qGDenjtUy2M4NwdolSY2z2oAzLHHVE4ydW8w0whokXkTetz09tknqZ6jusqH9JSZZJb4DnnK
Q35ZCjCZP3EUeYc96uIa2IRbmXeDSGydhueCX6VqYctZacHVcJu+qtJRmU09IxGKyeV9uCwCP5uP
bCeOcdrlN3rWCZfXfrN3TpFMxtu52Q7mnSI0k5EIX0ZSwa6oD5Ru6v0DHMtuXlE4NZiVTghaKbhH
9jEuxWIT2h/V/9JosnoquWNYPXJWLdcFNucEHeckvcvYdvb4YRYMES4nzIH7RgJsfKKhGxY68XFZ
vo9m5tGd/ltXbx5qHM318sFDm22LbMseegbcFAEK5t5ekZGS38t51xee8UPaQ5a+S82MeeoZnUWn
Ydck5H5V1xhkMVjg8vQcK36XIc52Zv1HUVlomgBS1TtzW8axmmPTt1AfSv8E4dcUTOK+g9HryFdR
Hc2PGgkEfMrG619sA76XuSNNiFbE9v1phWZvOioGb38TlItrkYRRCT171v3ALekMsrZfvyusJU7Z
IalCFS52hVxVi/T0pcxbXYigFwjZdHUz30EraQdYGsWroMVqZsI9qoKjVLdCxexJwog5yi8KuITl
tjU1ZYc0/qMkNh7NZDUchCs3k9P0lIpFknd4cdONqmVxHfQWEiRTR7wjnpVTirw3JK//bYdgTuqB
UnNt7ALNDF/MN0EjIJ5jLqKTY7PJT9IDtbhTkhR3q1cfZxV5TGxOuIUrKxirYPVe3d4/iyCOe2/x
d5krgeIvSsuw+uKRilOLOenNNJRjJrbmic74vXm9SyqF9zZh/1wpnoup4oaVP+RtZk913aHaUJcU
2B2ySXxlR7gP4gkC4gVsOqgvdee2CiQCxCo5tUJs60ZW49IvuLBXtE9wjWA2jZNdYuvXkwJJikif
wCcsNLwOFgEsC42mmB0CDQoj2sAGEvuHQQT1dg1/wuYeyTRg39hNXwz8+Fft0nwlTtZ9+cod1Bv9
/U9VymqLrY2+nkXArP/uknstGkhOudYCDQBuQNjjlqZUY8zc6e/QzXDFOAhHUv1LzuEdEVQSgc0m
HZFW2bdylfGPHBCFf4AG98iUXL714sDZUWesB2nAvnZk6Bjl0a9rYASRqJGjjjBd5uyuOoJHqNde
hEOjbrAbJrTUOqCSIUr/lbAiPlYVGl/ExqZjSnmPUemMSgwWYwVlTxq7+gHT/CNH3sPKbyRZPDbt
0ePC7lRPrMQlMkBg14nERnAUKG3kSMEie2b+86M1qFD79MwxrNgb1I38FIJZLBu2vaYhquS1wPIs
Lh7hnvFvNU+Gfa9iBNe1PjN7NjDlqpMs3T7j2DXcwRbQiFiG3C3szMJa6x/E9z7D9BYy+oub1o50
7UPIEa5GxlzjO0WMvFMOIIgx24q43wvLVbeFY37AR3biXWaEgtvJwRclZAYe/mXy0ZwEn5Ao/9nh
w1UyERedF+2HGw2EN9heVjDAEtPwHH48jd2VAABVXPDdS69025d1+swrfk9nMPz3/vovNaM+5ClX
Bq/etk72jxaPMUGPrzLPrAZ70hK55Nwx/xcI3bQvAPEInUnq6DBia8tmPNMdRRcu47VQf9LZ8T6s
wLHelI8J8Jk77v6qQZBcr6eKA06LsIf97snC4N3uV94Uw/EzlygG9LCDeHXHmQxLoJeThrVYtVfp
zaIJ8nQPbWsnU9n60f9b7Ylae6BuGsveyBckLzkS9ZMTIqbNKNOQQm8ZP2avWTyz5RbFdp1NpiLW
evNXFnUfUGixPDnjq/hfk3bptdKeKMFAgY7osKSef/OQAllVwkjl2YpyxwXsDKdpOd7sjA+w8nyH
tLPGUpynHCkbQSbzouKXQ4aPeustgNh4zhv415GnMN526nhYjgkChV39ed8nJFSiriT11UhF5qLo
YWC1FAv060RfMXD1oTyzU0u/GFasY310Gf3JkFaIRzSZz3qYBelNzDg4fAOV2H8EOPShhCF6TBSe
Po6KshGgmrZvBzAd7LaWlA/e36O0Tx+qmRFUAn+3rUAPWaqK7W4m245JkU5rcGKfBiXy9l4wAwfV
j2VPYbT42T3sdPzGDVSTqHDG/5sIsXu0e6iX399FSmO1xZLg02qzZJsBgUNTMmhaTZIT7kU5JVRQ
1nQsdThazRIpYcKfymt7DKLrLoogcaVXYME3YN+HtWA4Zb5v2e/9SWkeDGmnhDeKwNKwxvxauMdC
VBr2WnZIrudwjEAyd9urclxnUk1A08DsvSg0PJg0DHTwpvCHGODdYNQeB30csQzrrU+brpV16QXG
7BxQyElMs4/oK0sccJXa0nbY0hkuZofbWnhyXUmk0ptrJVIUYYerk+Q3eJCoT1P5V42/7nWixy70
zUlMlcyWFrC/Z7d674RgHWo33XOotrffKM5enzqDrY81ogt6CSFQ4nJwpw120f21EZUwCENfWL+P
gLhOqyeLKIcI4qnfg17dIAqw+ZX0qtaFyhBMlziHDIsq5HWJYDhQLw4+OKxnkQnU0Z4QOtMmcaV8
23kR5mkK3A9gwIchkAI2d6ytiQddOnchiqCueUqgjrv+FGYmAcEIM0kOJBijwMqfVlm/K6tGHwJD
wKCNq4MYht01+Sy1nwSjyOjwP7wgAeQNOMUAevEVgvL+v0TtdS44NBqKehTIWPISpVVIzo5F/Ugk
95I3vX/DhJd013jOySAmGb1JLKs4YzCRXGW7+0TOnzjodi0tAUkg8GfDUy13cMac5pvYnq2A9XVD
YmbEuc+XPMiBr7AZHjegiv64oyiBkRNfKkL79HLKo04nqZUsg6i+XRkm03MLgzUEW0Uzjyt9VhLr
N7deJPFbgH9tsl70r4glHL4IBb/m/eDaizJciLlE9gXdGre62sY3z7RAdHUMtmesNKhxVXSDhIZx
FGMhxrUlMCx+sMmVsjZ/+8k/B80nJoeKefCvL5r1q11ZxZxIVJdxpFG+DlpjB669vfW1DrVftEeV
K7guqm99XU9pqt8Cx+WL2rfOUZhBoKbuhNkOaz/H3aps1b3C/HwMR3Em3gv9pKUlKJoAF4hafSej
3zGq/zgk2zcettDcT8/c5mENyGhcnVnjcUESvRlAaG2nLVEqirez8J2QjVWf2YV+4YUA5rElg33w
H2Z/3KyP5qznkidJn7AkXiYBjY7AvOfr9YvUE88zfi6epY/mKRoUTthlQMrxPTmNkuCQwwo/IHXK
Lnv4UI3/AWLy+3qNNK7r+xGNi/6fcTPucxIhnph2eAiX8vmHiUSq7mqyTXMg6b7desiY9pker3++
stvpARoXphSR0aqQU3ettdTPJs5EWyoMJ947lUiQKdnj2BgM0W1IhIzbqsFcW65E1CbNiW+4+3Gi
NqfXJ5fSUlGjAKsDE8wInzFtVH6yQFyDLr5LerKxviwDbEfy/RkYZQTRPupEn/gQPuIRjMSQnjRL
igLG13qbpE5Lwx2TsPnHUYyrSHEVRnMkp/vCtrGY2z8MaTmoOuGuEY7vSaDEiiNquqlLwIwH1gAp
RSb50xutxJ6NrJWf4S8LwoqXwmkp/9EpL/DedvkCcw9iyw/nt0ftrBRT3WnWGsf7I9tgeH7gR8Zq
5HPCjSCrcskbGX6bF0STay4Obwh35310+jcPgIgWcto4jZj9QCV4G9h3q/XQVODrMnlQ/zy9lca5
FCrqGQIdCp0VOs2a2iyl+BwVCEvcInILlitzn2mCTjD+hlAIEGGr6TyWwdwtOZo9rhVqQq1wDfKt
dRWFLiwcN6eR8AXuJJh8cYPOtI+JAWVZjCPVd6tXAaO222dhc8ExUBPiIuAbTVRtS44vQ5Gu6dko
zcOQK8awqhkBK7nMg3QKw7g+91H6KXG1CN3Id+0xnORF7E3MDyLBJ+b1RiiGkfJNQnAzBnaxGuRI
eQRDQNCRc5NKxngWmKgmArcfSvEzwAopRLlYtX4TQVYqKbIPE+5RUM/Zj40R2rSq+QqcuA3kXhle
OteEmRZnF7IlKHUzH0TMHugMLFudFr8mSt8PNJQrsW8sUEJPvN2ND68zmoFcB8pZGzrfD1UMoVHN
Ou6+mIcWDV1uPShbPOtodjPMlmUJyy5V/ozlSiCqBWVKi1y4Amtm+2xzGeuTUMkgXpAG9tpd1YNq
XDTSuOQP5AfA8eOoVYFBIwcZ/tL/gnmIKtOLICZWfbtVY4vGy8li/5Z1ov/2hbgcHllcZBQh8xcN
O33yecodDghIOjU80eG/YRWJcYycGyxC94IvEbpwW1Fqdd9qiI67pB6944ru1q/FvAtS27XKq71L
/eHqRb45bHm4nQODFJ1GsxXQ+5UeOUK6MgIomnrycm104vghI+FZdm22svL6U9OcYJXtDuSd6aTi
YN5kZttLsfXkwgXF8YRjhuV0R5jAO7qZoOp3a8u2aR4iunm7stPTMkCGw4qXOtCxkGbk3K2vcXwb
xaswgo58fx2nyadvGp1AYIB9s2MGIqmMEyhSc022HMI8eBlweObPnT+yM+Y7IgY/dEGM2s9xcx1H
rocMYWjb055rOyg8eTO+jRyLulm+zXm1QRGrsHJ0wwh3zi7MMhgEEETOWw7KgMixksUrvtsoY3bU
fIbDUYNHtmxDaZOSvNBnl/QhibxabDfFVe/SelUe2+xsxwPjj3ia3kd7eiW7HHYgUe/JKowB8MNx
8ICHbdXQEqoSybhN9j7+L756/D10LQGpVWonJ64psHQTaN2MOLg+oaztVbe3sGotTYECUF2SxbU3
atlOasN7PjO/ewOKVmb3opoSlOYNgxCtDmerGqLhxhyT65HqaoNoFvtWYR3SBuBTPrkN/emlcA0f
JrQ3ufcvQVXCr7knHR2u2XEHDgbxwp+SmufnRDaYQRDPOwKjQY32TDvMOEGlzUH/lXDAi2a9hhLM
rTcbcpN3vxw2wiBJfJvUG16yjshySuAQw1YdbuNzyjvNcYEQVDZVNpklIY4QTbGgLnFyDrn57KH5
ffX0MozaKvCfTyI4mDb+GEWZYJher/gY2lwUTh/AQKBmUMEq95548KVzwIPuvwIO4uzz4/bf74yG
PK8Ms1c44D3qTLk22elNRDeEULOZ3hcyMp1bJg4MsOTiluQ3ZAc2UmajeQdlGNut9QJvmXA/nTV5
5WHIM/IYfCguCF04YKT39JVc8qy3NSrOoz0jj7MI37GFFQ4IRyocgAhlNmwk8w9uhT1n5BCXCOOS
AS3hYxe2cKzxz4KbmPW2K9Y/M8FR4tFod/b74tOwWYhcDnYQT1q2a0+BuSwiI4EG6TNUEFYSEqVM
RXILLxTf0JHG7K2AXhV+WIfS9Vl0XrREYP3q3/Zq1KSZfJdVrgcXyF+9BFDam/iPwWd8WcTb0HeC
MJYERfOJ4NYm+C6adiqB9UGliJJtyu7m/KK5mViID2ZrbzcwJYRpNEY6n7XxM/uvWKBEUDGzmNDe
58V1YNEGIBwV9Dt22pyiHAWONxoAVS6EOSryOzgI4NQqK9HOR5KhPmyQ84PDAkNkbCF6YTseqLpA
/sBsWltzTAXiPHUpJE4akmvlmuv91EKdTcrPp8Ut5N6RszN6Yj9was9/pb4uQKaYXjqaSypnQy+R
j5UkSc2H35tzFviREdbRcZ0zujzZtb/9Chl7KAqjtgft7WBArC2kMRLdb75kOKHrtaM3Qyg/uHeD
uKroitAp1ZiVOccLeNIatMcqfSUP7XtKExOFvcvqNFHEBxxTx+PnHEJMSC/uNrpdnK0aZ1vaNUqc
V3yJvfs1Q4pPuW9avKxtau2Ie83xdh0DAgzYUMW4oqBc7FHvyl9u0UIeO24RMHndC726eqQknCrk
gvOWqalTC8wyDOEI78ICTinNTLFobWcRqLwGrhYvRC3vx9oRpMLn/XBAgSvnbEH2w4QT3lAjxvDT
1VNAA2twossv9vK5COyeiJ2J7KONCKgFOyGMS19SoXLgp0QysUTJIjTQXB7xKnDGsi13mBT37Idi
uHoaludfnTrVXRpLnJXjUEtcjEWIumRDBiWOB2AuIGejBbLq/8SpA+uftUdclKG0UoCYGKK6K2RY
Qd3FFzxDDv6JNLOL6h0AYF5B/rCLbG7lDQXw9o6D/XpPBayjmWnuIkBboFbFc8bN4E9CJF18nLnh
+vLdTWFgxOFAmy81CSjKrZvRg0VIuGyFYB3pJShpSvW9Ekkoc4wOeFXSQwTNvAPpl6HdWZwHoK85
0cYMwInREITBm4GqmHSp2zhA14TBEi1oRSFyORUIh48KSL0L480+0ySkodilXA/oHQ58kn/mu8cS
KGPumDzEeQgq2Z1DB5/6jOGZXGIS7PkOLu87eMvZmGLDyM2sE7BwLcT/9P7wVXVJ2cvQT3E69EUf
gqWZ/w0Wxz1jd7ivzlsDiMYZjy5HmmzO2WXh6NmQAheZ/vy34yUotPwyl6CvcGqTQws4PDmbsV6e
MhTyjcWKrs6gde0FVPPE2kYporTpQVkrahEfPdwVmUccifmJnGpKmLb5oZv+5Z24aDyo+m8LqM3f
Zg8rw6Y85QqKsK/jjTcV2LXyXSg6ZuyiqVZMTxQov0nRndJ/z1AvrQPW3HWaD2L7KcEANYajruN3
XM6++7lHFr7msDbSC5c/9MxKa5aHK+P5AXxzs5fnr/tPozNByICMyso+/7fn1v4HLqTdhexBWNZa
3g9oI5lTq4tPLvXGnAp1zEavNcJHZ9zrqvENwMgYIco3P9aVesLQQvFLff9dIThYvZGhxqHHAt9u
70HplCXUFGuMwB9ysly/NPOf4fqISKM7QUOVA/OyZHcyHXTn2GdU75RSy+SLoOMsXtgpOiakOVVM
FZw5N4hNPCOXGmemrQqWWektGGYcBs/vQSZyHchVf+Cd/hDIkxF9QlWKZbCRX/iYHYmTVWKkgUc2
7HVzKeGhbsVnpoFwcK7pBIR8q74wloQajtx2u7ebje9RVZgVaOJtDt8tyc5X5bk7uRIvxMCyWHUg
jDKScg4/Di6LGGMpG9VfA0PMhKv6QObQdUaxMU/Fqjn6pZVy/5hOcpcZ7Wqqp4prBhDq7byZ/+Il
KG+widAo0Qcls4VNVbF4M1Ct/mvmOIuz3s0s4odt1W3npokMw4UzkatXwvPfEdgS9LDvVfpGKmhF
rZvI6+6U9VM/wPhrnyrI+x2sv8v0K9sj/AMsKMIw9bh6XuqIq8IwRZtm3cQK9CyFJzz38K6pH4W9
Akvq8QBtq/ThU/ad1sOMpIPxVdD+sz0f5G0X/nCIYxd+U/PKztPwPIp3rtf0uK7CLD7KarMC6PKf
fFxXa3yqvxJfT39gHfoDfoQxVQ+ztHe4x7XHqzgq0fweY6xHZ6A+07+ayRBaK38WYnv0zM4yxGGj
ZQp7CZfbb5Vebc588zcZRa6kKHhYvQd6FwjMwxLQfZbj3fo5BFECJTmqo1HqnO4HRFLj/0/Jp7Zv
wk/eIjGPnVtbWB0s4kQ7ITDxf6mW0Rc/0hr/9GTQLXoE747jR2nwrhNgQ4wz1zC9jPjhf0TFMKss
kvQijHzSX1P0lnnJzxxyMr60aJiyjEBcodnts++e2Gw/TguVMh3tSTyam8m9/gZscoE7iFLzz9if
23UZsUrITfiraAoUDcr8kR8DFezUi2cxxI2QMrjqH+Be1EciyjYRE0Upg1jw7nkAEkblHSwg9F0w
Dx4vieIZ022LCgkOLEUnNJNPTHyRRfTuhOGt+KOOpFykJTDXYQc2cFeNAEjE1toBQVGXcyNEZK69
TZutfA27P50jowdDyGdTPZV8fPTLdLD7K7eZbrEuTlbFtz/h74vepzrv2wCfxyhOawIpOFemEAlb
o6U+30+1az7A4xM4e0oNl9xfg7eysJpdhJhjSQxGHAEmz2wWzAlXaJbyiQ0+VuaMWnvrA1h6prvr
HeJhD5NJUgk+QzRwE1YzHIhT10Vd1I7CauXCSstsn6mTTBH+ZDh18CgvE5eePOqGww0Eg4bP1hdJ
HF04Yl6Mn6BggBaRcr/pz3UJD6rZyM4H6Xb/7QdPznwODlxBhPh/WDA3645sZBBKhUd3sV/19oiy
gU7k7HcbKBRefv7Q9aOUJ0iXhxdMIajnkoq5IKhqL8ZQq1JbyXLYQzk8RSMyuyJr9TTOcFEOJHjD
rn14hCxhy+enhq3aTeb8RAwi69n/Oz/cPJgAgYYmTAijb28nviYT8SP927cgWGYZx5f1AuPZMq2o
j7yasq4aUCNKenciT+pVXcDrSSy3SBLaXb/MSy7Yu930gIBRg+73C7G1VvMUzKnunaydqjQRCWxp
9R+SYgvhnHDPLYqYWqsXnRtXlNVUTGAbXGHGkyD5ze060b4DP60tjB4j1ML2hWPyunbe5C2i7raQ
ruX4iYXz9ipXAkcCPqmV1heu5QozZ9pPDYwiDhmd0ubKDU7IcwlpIqD5O/pwedXjrjAF8HjXGJyS
C6GQn1Hmp+wkCVYvBY81LCN1E+186RDQtrFn+vAcF28O9ab398QbZIjAdk+GrkO96vM3SKQ8aHsP
IaRZp3k0Zx35qIJWV1ntPzQuD1w+8jGxh03qspePmpKtbRIaLI8R5N85Pb8W2Vv8xk6LXtx/x2Fe
llQe1CYUkGO6Q1LahIC1TSetitZD28gSeM8R3F7osvqV2y0uuJlOJ97I89Ql6g6NcDNVGQcRHl0x
NhDS1Z71PPqATzCvZjCkhMX9cT0jpF8PfqRVhyEMOodNmga88iFSHngpeHUe0GwWLMTfep6CddjR
66uObOXYlhF/IRh/TRr+ZwE/cklnyR7FYvDSSrQKnD6tWGHNcXb4ThUtpcsWSlLXCs/MIrJpucvk
B2fcopvO35xB3cj35NvRaVIhDDu77whnHfm46aMHdeov50Is+ADpPefA0p0OAGdvnggahtM6wBIl
PeWzljGgNR5aVfXWJUd1WT77GkTxjsVr4MibbqB2Y/MrleUfkCEWWsJF56tXkLp4cYHxMEqlP1aL
dm+rS8wnCiF8SullVaKlKE0k5lXt3NZwRAIGlplWz6MaCcDhnaGT/r0EFfLN+xq10xDVDsE++Pk0
zS20+GZAh9XVjJx0sjCSXdUVg8nK4wCrED0X4An1V1br1+UKHhazXsokgwUlEjtF9LLsWKdEGvqp
Z5dEHmYOn73o+zzbM0vQXcJYvcD+nMPMrWpM0YbF8KSCLocaTKEVJr+DAeCH7TtpGkgureePfnMM
JI8rtz01dRxFAxbxZUdnqbPwBgTVuqHYylt3VldbXuPsqDE+q5IuB1AU3olpzhdfiqDFMF3jF+iz
+TApQh9JfvlSO3LVUTzLwBay+b1F16cbs788IMAg0ouZhMd50tUVwN4xBQfd2HpkZhc7x3gTbu6j
5TpITtnWKlx5JHJEo9REXou7AVGWFj72sbWEUtUyYYq8fPTzDkZJ2vuQwjP59t0kBjDL6gs0tIZg
anWeVD2agXrLcALKLMk1Jv2PaRN1BL8MZI8i7BvN+PzSXKtkGvZO4tBM4VmLYoefC1zvwupP3Wec
nG99x1eIG68Q0AaIy1jfzzOy2ADetQQOcNSnt4PdXYSX6E3Apm4xx11m8AWw/SU9sU6nsk0cRllF
X/sL+4GERAvH+YwNf8v6Y8l0dhI3O18WrYyXqvsEPsRK6OrjiP3d4m59LpSGRzHyowJAuEv14jId
OL2bR2tRltrQ2PtKp1IChrz+LLbFNPv5zC7rmZzWDHu1MGt6J8BHhEbALoBMm+JgboNxB4FeJlKT
rI9wPjLVesM8V1ozYEW7w0ZtFUmKglcXBlTZobLkxvuXR8p/oQGQl97uykdPNawkG88/FxfxLKuK
rdgX0ubs7oVkD+vbFeYNM8eNwAVDOLztG73q0jVaSKp+hwlsHOgi39hqSekqJCRdvRzs2kJ8geUA
QgQGF+vkjLgQ8gb6EadnBQsJF6APmGDCp1NS6X7zw9PdB1NL1SscbGx/bP1K4G6UGLrVsCZdYqbk
sXV4iEp9bXoxwmbPcSDtoRB3P8LzKX9VjKErhTvL+71oOWgDsYo83CR6g+cZ8RHn35RfyeNk9ICO
EVWEk7vJX40250QO/2MBH8ej5FGodr76ka9cWracuEdKiLj2LOE3Gzf6RkP43mdThaEDQDRwHMm8
8O0rg/8roJIbL/CnUsP+OULD5yHQn1HF3XYPqlzEj4s/u1m7YT6gsLjQ+cO2vYUJ+YPq0JHPIvmN
S9RAbn8rkD59OYVDMhoz/Uah4R9OaVergIBNEzxm5OzPWL6ganXipOI7EPuusZ6Tn11GHKbNn2nt
tbCJbpbkj9xKz0ubNS2A/7CgtesSWrmeYXMoenPVPcEu1brzCDnPUbRzU0baMS4adrUfXTqHYpR/
A/oLQzaq42kNe3oRSFCrhRusVEDyeP+M36reSMGUHO6P6WJbBZ749/js1GIIuhfe+z/FC9rkxa47
GVRwDeIaouGL3ihdB3AbWOTpKh/UgnJXLAddQu3Xtyhx6eXSf8MrQN+6mw6dGOhYFuQNMKPVVEyk
9AkDGAZfFtQZbcyPZBtikiMj3BNu1t4BYhZ94NP1R3n01xfJxPn0PfbSFKLiBWr/RysukRk8MWut
8yc0HXNCegPn9/QiNrcQzVpX7gG3rn9w0NQhR5yG5oZZPL2RVG8O4WDQQM5nI9bpWE0SFvkEA/ZW
0ByI87ns2ORcEyuyN85v56AWkoPg5WoCJ+wiYH7PYpA+h4fLzaNxoCMA7cXO3mH293iyuLfcMxTg
/KCiQOwVbCJtGo5zPosk7PgthCqKONXMqLbbTc+cY03VwafoHaah4LI8JtcnLAnpbuaVxMZbY6Ui
Doe67qtqPJpdJuIQbEn0Ce6kl0D/Vw6Pgc8iTdL7i6LrN3TQc2YQsDyJlLqfcLptxegd4PEIkj1d
K22BAs0cfnlme8lvW2tDuzdfFQGxkyFHe2ONEmr/UF0MWsN5YB2Zwpf1vyYw9TEKsV8CQPib0mwJ
tGvpj7zEWMSMrCXZN4qedbzH9AvT8Gxk9kO+Vw/M3IHKXbtkoSrZJJc35tMw1gx2QItn7qDZ8vQf
yJCGmbOF/72cBlkgBCq+ItHAe+nnKnOngCi1rNcjpWw1tX3huaH22HJOmNbzLoIOEgYRhArqKa5U
cVbBOIP3aXlhDIhzpa+ddQU1B3Vy5AqP7hZEtQ7xYm9TL9zUcf4RWTuvTihpeIIsvnkYPZ2YXkkm
iWFyyqmfBMJT2k/mXoBeVfwaS4Hv9spbCT6w3BUu3267zG6QnfqdBlfcPOf7qLoH5mtcUQZ6pkGr
JnMqVOcnZITue7dJsxyuU/Edhtud0O6CHW8TURnX+MwFrLDb8vzgYFETUhWpX+VgsKBTTeGzG/tg
t7NKf2LIyAW6hDAwbio3P4qwVAtrKiNUtBkWmf6V8PZR8nuNcdWshRtXwCFk0yGoiwADpXi6dSOK
aKmAhGx+vWU4VA9gf55avXEsxO4ssVCfb2BA8ritP1MnQTab8SNqKtyu100hyN5UP71AMsq8Fgn2
aSAQ+e3uy7o+5mrYTMSBLrIvqh98whXvOc2C0AuCBbtCrx8pJPmvjKEZORksnxCus3+OO68OyHIr
fdFl7tyjUxNM7mDkDzz5ESOKNz/j968L61ZuYUw3Axmensz+MgT1VGYHDHyCSGYllQGgpWrJNIBs
NNt9TVILPtWjKd0FvNoFwK/5KBRNc/qND67eGZF1a7oE7nBzPrWI83V3xLpCyPadEDVBVMaVNA/Q
2e7X6RaaYPHgQa4Zb2WqQrLVNc4QcRSXHuJtS/5r4F7jWsKRu0jg/wxLIhj6WidEIFaLrKwnEzpP
Ok+7BdAf0jHY/AlSgxejY//zRPtdKfX7qwIg1N6z1Pt+yf2g+qKWwwvGstEMevow07l54rvfri9L
gRnBuAjLkMnAnsmJvq0AhQyhD1rf01SrFPWVoXf2Or7tfUGPsIKTLeRUwR+inO1NXFsTTzneIxZx
jMS1NZp05N+1DwXt1fzlh6lXZ3RpCfzBDzw7muDh98BRyg8teRcgXO2zw3lES2ZDotUHFbIyKsEL
+buQ6MsUU/oI38whEQ9cRYh9+lxPpdaSLP3ms2J9P1uDvWbhGQckk4Zpc00tLykbTdGWcvMMe85/
8jBy/jAaxuW3xRAjM5LKS51sfMTQog/1Ce5mC3XlflkdT6tMtA9HQffm3HzndJDlK+msqPFMopno
sUNwyjy4B+1UHOSp77vML1X0yRhpweyybRFzbO72wjvm0Zu/Woamln+iw1o3t7unXYJrklPXb1bh
116n4hOYjEaY8xDHCuvldo0voevikuiCnbZEtlxMIrIVw1YvZZlvrdWj2PA3TDstesU3cUQLYqII
r7HNVSmnKbty6yHwsgc3E7hzg381YVxWzHNh7p9gZ/a4Ab4HQfdsKcLA/ZHz1HVebBqx77BNeCge
FE8FPnZ4Tpecvd1ahlItYe88akDygM7bI9h7S8Y1ZMGLWJPA/swIkmhBL4mOLhiiAtpc7sOZ5yco
A8DDNE1v67Pb7KNKbQ5RLe2rRzMIOovvBM/ykmHrhQJpsE6fDxTD0nUQVPhp6U0xEv7MBrwUCAB7
yt6cMs0L8UW2OXCtS0q7fDt/YHMlUFCG8raGw03wVbZ7XWoaFTmXh6tQUKPPb6FtvYLfIxb8h7XB
BIEE9ZVlfEUedT0UiDAVFIbKfqmum9vdYLxiGxXFkMQv700tY4E3aDbyZTO5d2Mknd313fWy+5ec
3wapfaL1ETX5CvsnMpdsLEab755y6eBESaFYW0DhBJDXYImOm7DdJiqBqJSZoQk+WeO3rfHsXBsc
chLXFuQhw6sJEFFbR/tdd0iz2wNnyY5/daVovlq3Vet2DbnReVfWg9C/kyclOCjQJeVmTL9Gjigh
JJIH/esAIKALungQRyZd2YgIV0moiweb/JPe2V8ldfTwSu2L5K82az+CNrjwxX569RESbGOb05gz
G5U2xQLKFGhJ7oL0U51v6NMv7lUUdteE4I/jj89K6o/ZDmvdhMsbIatN8FBJ0Waw8Ul6h+Z+/tj1
Lg9J3413r39Ky4sOBUYpjvh5ArqKt5gGVvX9WBndU1y9mtlQWXdHtH4GvVdKFl2Iom5BGEVLLQTV
rHV+q3Vom0UX4t2NFAy+8D2sdYMs+4N0jp9GuFkvhHfPpK5LSULkKwuvOupBsd2bnk4DliOZQ/Ii
x0AoL3KylSyD8f7rD4hJCBcLDqoOdm6ffatLmXtm//bVP5F9gt9cUpOrtVZK5iB2uE1em+UYRyFf
deEa6DX+GFY7VLwociQv4sPrQ1UPvSYoExfDcH+dGXUZN1Yjs2qC+mKxBzI2bTuvrFCd2XWnsPrp
HnoCu8OexlZfkII5XxFM3fy0LIUb1n6Gg+pSF5ke9Ngx1KM28dWUMlzSSpFQG3egqubTqI2y06rH
Q5cXH/dCMZ6eFgMOVVpobGwa6OyOuLe5pe0Q8DvMVaoAcPMITGdJhrDXguNHUj3/NWdZmahvVtkd
+leW+g5Eav9707VHHZDubN+nDEh1xfnDGLdUIixWov8552P0rfb10KRCMkkDEk6bEDIec7kjgo5R
CHQH2GVMLjN6EwAalNHqtOWke9ceQGWmKhtVXPaPRqNfffUnUrH/MQdhRxZyM1bUIPz4MiN3hyhG
JNp6t10EAYrIQIDUDZGDyj0+xwBRYxePWycaoy8BBPfe8aj3GkcwMfjKHRjT04w60kXRPKcaibQP
R+OLbv9+saSKj3gQ+jC3KOq9Yfkxdpu1f3gaGHmiY9Pb2mqYLAMcdMzwWaer2uXE0dQT3fnEfH2B
ZeXyNFhfS/kaWZaszSijHhbOb4QkVTHws+NgvXd7tfXrJB9Y4gOcmybm6QpwA3yJSBI8rtyS6l2K
oNgNkOLfSnkNYJKLUviTGMpvGPGgljdzZQtcApPmKiPrviJ9qRivjty8mmBmngbXpbl9upg6qB0X
ySdsSUUNBMhHnmRcCTyHVZb18WnUcH8wixC8V83ANZ+/+hfgY73dPLec33Jz4GfjcZgH5YbknIHR
kXrRmi1cPL2gxyZrzSc7ofPoxt6hkv2/ZRL4fZbQEzSOe5emjliaCnW8bn4CptgEej/MzWckiKzo
VRim2ZNo9/cGCI2dlO97F3SZUTQr1PtvjjpbTi4bZAxlNqZeyI/vf61f09H8tlNEvNF1jL2MzdyS
0U6eg/C8/+NYnffw3KZKsOQafN3zssHAffcwgyd/5lrlPf0p+S6RAs8tL3LSdklWcHlsJZBMVOxo
9nj1pbpwKl2ksgJlsiPQXNrV4qAJhnqIl1oL7JGOcKfYxZ+ttG4nG94ELqOW8xmp7/LRPbv35SB7
71OxYFrgo8nqQ1i3F9q1aThPDxfRDl9ZQFNDGXUo0SzipkUg97dB+LVTgtAITGvzV9R502mkb9K7
UPC1Gqp4DGoDL2rXTkqOEPy2JB5bnp7Omm8yPZuLfU007zng4mq5GrsalenE1NmITxPjwVj94yQo
yEijuuPKqTV9K5BgHZqMy5M8NMbzWkE5okSQxJETl5yW8/GIXQhh2kZIu+JUWKUBoQlY5iWpJtTh
IWLGhAx+/1AvKKnL7aCGg5JaFlNhIQv5ObFzKZwAmhCF4oOAh0QmXPgXmHb3iaOMA8C9wsfUK9eO
p1+dClMnwvYZACabU0mEQwdEQH6+zIHmi8VmHangxlTywqi7GbIn2TXtQq2TrQrIn4+1rTceo9Ck
Wl+poxPuIm0/n1YqTKwWJa3ornkkChP2jgIWfTm2zyXjk7OzqlRlZ5FOYoAOYaMd/t82FFa4Q8Ks
dv8kfL0f1Vu17iLJ2g6/eeVXP56BnDQwLQAVkQ4xYv7hWXs9mgmtbHSnj+/vFn3SzXDZUxy3yVJn
bJr7rGQUWdfcQU1rjFtiGStxWMLSqOfsmKc1FF4rwGnkRb2jt5u2u+Z6INJTgrr3I54/TEnY/rqk
PkLdakMHJbvePwpqkZVi8vpb9AdCzftxkdSOV2ffxDDRJIAaIOxGrNixWT883lG8EGliZCHyujj9
fh8PLGHNsGm9iQRYcp+JbL8zKT9OKhUFq7ZpQ/7EszwjV0V5AuZgG83mJftbqONcctSj9XzHlnVp
1RqxK7o9ptNHFDZ0YqQeEml3u7mYGs2ntA3Kpipsr82w7NUiQgXkRWn/zelVVLI4G1vYzt3+6bRG
ontecPXdGsBge+9eZTCdI5l+iHcYxkTe5hvor0VBF2134gU2uDlJfS6s7cXxxWd2G9PBrR0Ax/BY
JZ7EqprPfrqj6TGXe85uXPoe6r3Dpl2SVhVbOY6KdNNAoz9sXx+6F48YNUg7LWIDovlFCCLihljf
34T0k3TYAuhFpw15qw8QCcYBHrDesGIMiG+A3r2O3k3wzPyaQARk+luR9lucwvOt4K+GvduXMCGG
bQpZXD7i1bjvxWSSLMELzOWHVU1c8IVAiTlHPyauWQE+BBZfJp5zbW1B8XsedeYRQ74djd0Hq91j
gppP7LToXUgG9G4Rz+kjNAy3nJH6R5mBuAEC7J3Vjf0rBdA1u7Yntf0KJlqsGSp77GvKcPk/y6Lu
5ZcN1Kzk6+WciAGWwzBr2Xn55tub/sLtr8GqQd5susOg5UAXhjLySFY2ioJgrIAkpc35rlzEappj
6ACfauP4CIpSVTYkoBijxVG0S/+pRvtJ3i6qF9IpcvdVEM9864VH74fsUwKvjNvVXxKLbBYG9jlU
w3cqOz/Gaq2Oapf0IQ764rHSNKd00uOVmReeTOuBnYa7DPbtTtUCyFlzdNjSuimWN4fecOpqFQKu
H2L9H0B2Wf+mY1/ibA8aSKD6CtV3tkUkRKxMwGxwo7/8RxuoliCUCuIIP7m9jc6TD0zW5CdfWQTt
EKedB85NGeX7m9td9weRcFeUQ/lnGlxesjPk3wdGZhEdbqx3OjjdKLm1S47k/sBCKTGy4QXzvkDU
/M3C8JWw7P4WYvOl2knPwITShS7mBwo/Va4VlWW1sJHb6OWbDuoOYZJJCkMbKLmO3fQ1Ye6N5GBw
HLYXuf05eEYv4D4Td5pDyeOpS3VD0/qgvajxVI4zivww+WZN4xFdBLW+uCnntN2inaKy8GhOKvOb
p7cd53BSqSGzBMeQgm2xk9GJ5IKNKyKDDVqdGMtil+9Le0vtMnTVzeKMg0LXTKzdRU3pjmPl3EAc
lvE1u8Ba+hbbWUe0lPshJdjWbufYHsRC92PZLGYZLNImbG2kR4ADOU5JXgt3oW/LQBh++bZUOnQp
Z0AEfTs6sGTG+k4ycGVL9toK28ReoxIDiXygYY24XWGkIv3EoeYbFuPZGpSQjfrQSLIWGTkDuFWU
HFRd8abNki4uzV3py5VxYnC1UYLgFnKUWGQmr2dMu1rZeE19aaS0H+8ZTJzOkUXvs2xnY5o1hua9
hhKO01ufMJz2ZQjku32M1RK2oRji1tCC1lx1+xDmxKQnvqPUoykB6ilHxtecYdGMh1r+gMFqD5p9
4G+oWHHrN+WrREQrdh47vBUl/otiFtuoLEWzduhukG0TGNKcwMmBPv3DmRZ8QcvBBGKG6IHRYLXJ
MvB1phxB5ZyHB6aXroNpvpKoPhuDZWDeY1ZgYwJ8AkN5U64fGte5ShTgh0RjP4dJEl1tTBrZolXU
UP2s+k3KBbdWaeysKZz3cbSXfd+/Lt1Ra0D1+kjhCTa3iiJ82XP2ch6IowXma5j7lT6DdQwpwn2Q
agiTCh2jxLhSpTJAR5Ll6XdKMqv9j2a2YhAI8hpG+cTxnUb7nSEp6tHLdPyCiR3KLR3fDrVRh/R0
cbOVQ8aukXwoUcBHl5SgNMASwKSDVO3ZRske5+3jwySzQZH+YKD2SB+Sc5/YuEm158Acv2QFIPmo
Xzu5T+DfPluvAhbmPJVLQwy8CbMFh4X72J+m8k1dB+ozw/zxQA6Dg+vHcIdZ3Ed0hjNPtD4cjHvi
BW6psqSHABxgfLfIKHSvO3AeP0dD2Ma6Pu3yOmXN2lUWJDBgv1uJUFHcwXxjlQqQ7kxDCx1qVbWZ
Q/BIeLs6Ffd/ufVqBDgPUvhtrhemfH/fQiBHwwNw3RT8E16xKNa1DfPz8MNjubx8H5mWvoddJY9Y
64SDJv/9NMEP3IG2j74gSPtFgqr3yI70CQe23ASg3FRQuvuNP0ArBs6vGXhjIR7y/Tg58ZT3AAJQ
rD6H10POPIbWBC8fd1jsceTod7DhV5fas9+AXn01yiECkfutA5bLQBbf4xLweu07mSQVtLNciv5W
xcGUz038xB/MaRq4HHIdtcQ4KFRGl6EFxBbQAKP38bxFbP/k9dzwSWKhIg47FGu3Zh7OI38AN1Xv
tuHm/IaDwSuhpwfTO8uj5VVOKzIFlgmJx3oVEpoLzqYt+NsMsx3WSkxcx/+p6COobMxF/Ym9g1Rw
15/6e8HAfj10YNmA5PcdFNv7nsgNEaWmUXX081WnBO1/eK7wcMuW7Mf4+5d1puACkFLuE/WOuTKi
QX7RLIgobuh/GuYYkL22rQRNk1H4MxCBPjpLaxkWzjQUNZ5rgn44+R0zk7DKRNYLMXMxEE/sHxG4
AiTFS078tL1XmA/AjpNp59si0ttEHIZhR+6Ow3qWL917nb5tYN6ZrQ9yu6EQqzl9zP7mZfKbLFPF
yLdDFOfWE4AjJycxM2HF2wbNE0gVDYmcBrX16oV46w2HAKQ+a8zStwCOZqsrG0kNmtAaU5a5Dbas
RQC/hIq7GjvlPUzSBs6LP//y7jantPCtY5k/Zqh289bB1mj1pFFg9kf15RagahGtqYD8Yd8922SL
4GSTklig3QWU3ZDUB+AOcOd734RN+NrRPhuQyFfn4oupO5a4ebkqjA6pXwpuCt/W7PkyzQb/dGKU
biYbLTHGn9Vtj+SuIPcBp21ght5mV81vpFEOMifKflAHGF7E4mzLdlGQT0jPEpLBvtxnTU7Ck6/Q
b7vg8tVgN32Z9SMtgUDOCMuNN7bew+1why4a7C/0OHgoIbfYU1SJhTJF4wyiMRcFoZNrnSEwwBV3
D+ylTe3nJwM9W8DVbgOZbnTDqXFtWLxmPG+3X9rltCdL/2KA2Y66U/aOBuOFBjomm9kyo0y9bTQx
pQMkYiVEuz1vzpyOGz92ELLJvSRIpLImem/gVR+e12/JT5iaaBqe6/H9tzeLNQpA9+qInwi5jCHp
QBSkBs2PzJ1PeYGXZM0XHzUw20YP/KGROKcxksPxlVr2UmQw/pIF8WhAzy6ue5lf2eMdTDST4/cz
4TjB9tJa7mTC0PsYfYUA1lft5P73hm3JSATiBtQRmxjod8rqpJRnfA444azP77Kqh+Jl6ISVszSL
4ur4zAL7RHNSkV4QYKOhQRzeivCNJdTsYSpoYjmyaCDc1m0NCIOPYHPnMwdzF1+FPRSm0H94E9Rv
3OFY7GMqVbpuvKMjRK1gD/m3RS1XRDzCiHM+D/Hvr0+b/oFGqV2e/V7DlwFnd49881Q7h1oi2XDD
I4O5NzqWyYezrTKO5dNLu8+Sqf+bZafC9NxTARwdGzmiTLZ6Ig9eg4ytvT8BBH61BdnyF3vAyfOI
ZMU6h9maKNRFLehE1qWG6rxibYzt04rzZbIaPwmD6eOiqVp8z4Vz2d0M0LbMWBT6vLUROW+vRDoo
jYmruRK9kRi9YekbxdsiCMO2EoIp0H93qJJ0dd7O+LcnKWASio9aTHQmxIx9iST7shk/tXtz9923
BQ9Juf7G15/j0UV6qFnLQ+4haXTB5BtT+sTJVQMDrg90t3acO1rI206njsETQbhuIcLVJA7VFhXg
Q8bnoXrUMq0kf8BLBpoZfsyMVrAv0NH/7OCFOolusrRjMqfLilz/YjIu3aHeNokj2pFebX7EWLHP
uLDmsPbdzhcwnbZ6EKyfctSrq5g2LwH/3pcL9jdXiepLmALzbPhWxspl9s5m8zSrJ+UiLwkpWQD1
2dsvnaRuNh5xLqnU1soZSkxh4T34aqZbklzbrlbtK/NSgD/rggzgpJonHuYzAvtsQifYGZTdA31i
By1Z1Pv9c8xTpYHomcxJ3ZPDibLwAmlW4TTv3KDO3IJ8QkzjqQ9hwJDkql2Rn3d2XXsjgm78cKG4
BHy8IzQ9guopZiaKxGlQTm02k3wNMFq5DWGeTJaCFjqvKEh1tKpGmCkMc6fWOx8IStVecMJZvSGA
r6R37UdY085LI1+yBgYK5CLzLlZPZlE8h6rxRjd4mR+QD7O07H0uMUHbkbLcIHjrpSe0SfUQCiBj
dFr+5Wg3ibxoTzPOO+MpX2dIPfyypMzOUUhZ4y7+oAfdMch+A/5dAPJ1r558v0yp0vPaDX8UMJHG
6LkQ3FZlFZBroz6RelHu71y1nIDlK38EqZ4O18OMvYVlPUp9F86S/5wLTcXPM+dkjI8cYkefmUGo
E4rKc2BwznIdfLx9mVaDdgIWHg+SMajU8lVJX4Rod5Z8OjA8Qx0mfqJvq6YQAAsG73lMCPd0RCxa
EFTT4QdsefjeeoRrpLskFndMCBcaXqT5P/PcR50VbJGTWrDlzDPubocj7QnmQ4UU5zCduhv4KHww
wLkzbfAhxNGGvsvhxBDqcyfNcs0cDBMCmWbzMtgJZIbinuVUysrqqQq+LV7xJ8BprJKNMrhyjzW+
dF9BDMf3L0ry84UOQ8Po6pSWL1xo4Kf96u4+O67RDHPcTBU5r9H5WKXXRvb3sFBYqyFPfcfnwN1Y
xRyh4Gfg58y0fJcxK1QFw2kUpe5bHGxKl+xpmRjOhpgUaKIQvlwG+M5JOHnUqudFGsQi2/qY+T4/
tcsEpIx9wu87aae4AKmCYqb1gu3y4Qbl7AmfivcNAyzNX86dBNLa3zwrl9q4NayLCkVZ8VFqRAV7
Avpa6wGeDkvaDvc39AaD3O0rR3J9Am6ZVTyQ3LfAQIqjd/0kQNAcjHrn5C2pmK1Fc2ewCuZmMCD5
iH2N4R3XKkjClfvBYDiOmSWxqv534VQTRwmKf5KizVsPUbC+KMRgcqkWxoFPEd7RcRXW5QOWRoOM
8NADvFojx9h76ePATJQSRWr2ZsGsGWYl7mjcvnDqN0yHQEvGzX62yC/1rzK8EI+GcdoA+nGEO5CP
Z8Xl03D6LjJWAJdCg/bUmReTV36Syd2iDkERKL0NwCEWF/z9SAh1lwEd/fQzHLQeHuHBJz9GJSUp
+9MUEH32l2giOot1rtIYZsNS558bu6/Rb0/a1AoaIJT8+e4oy+zTGnOyZ4cyBmOd5S/RkMNSMyd1
PMYQuH/vdIjHwzN1R5XVAIUZJo42OLuH6z9aId10h2g360Q1qdyDg1x/0MNDg7UbI2AMoY7QgTnE
yqIPDK+fBDtRfiTPMamjk+K5CGuPHQL8WKtC/fPSaWI+u9Z/Ubuxpznhi3eeh3HEU+YpUCCOxa3M
cyobF/ziSBm0Wve6oNKj2lf9pPUvtoATJHUl2HNYRqVTLsN+3byQf+3gBo7Woyd2v5LCnQ6Sjw4M
8ONuV6vU0O6b+7Ilv7foLPjovq0IOevd8MLJPwrU5Z6lOBBDvyFM591Y3dQHEokD6AZe6ynYJ3eg
qfZ0O8yZZiGAmFegxkIfr7haGIV+LLYolF18s2hNyv+bmg/zKnClJVVoSE9FIpnLSu7ORl4PyqeH
pTwVumks2bM23cAUMN/mwM3j8fPNZtdrBrxm2765U75UXALl3pREfQD5OH96gVzWhK6YE/1dWzXg
Yr4aGNbSEEFr02vrdSMYo7O8CXfmzuuVqqiXd/51d7H/1N+Xc0vgW9a/G6Unw3CPTlz2LX+HSvj/
uxRrjp4rd8v6/sd5IK4GpvCshcpSjroR+ccLShKh6r+4KFA+ElRTuV6wNnkHe0ytynMMlD/ZCGcY
eMP6MlfXSFwhaEVWUFflV5SKmCqCfBmqkidXz+vBDgN2kVwERWIXy77Rga1bFt8BpsEtZy5STyhh
7sG3X7rQ+OgW8prTo/FF/NsBcBiFmS3GVi04iCEIx51+Osinmvb/5S2GjfZ5LRMDLeJ4pNT0NNlW
tcDZornEADQoF3xsSUy3AVHLpD87TRJmVrwR+22C6dHlAer3v3BupyCwcyPrc+mRClVf3S5wCDNG
ivqRgO6+ZPmc8+/xKTe3mhLItIn8HO2gVuUbp+GW3FK8F2w7T3+ncVhXo+6UiRTecCYbe9k3W942
2li4t2KJvNOd3xTv1HPQSjb/7E9w7iPuP56ZK0GBSFXw07R1UMPnM6f6/p/TNvaUlUPJBzpr3XjR
IkvacxPddjuGUEdRuF9uwvGYqTrj6byJTVJMbdZ8eCJPmh439rbLLchlya8MJgghDXevQcLTMDuZ
9nuOkYKk23QZ5s/MfaCdVcTTWnmBeFhrsYU6gTm2XP6ta3Ef6622MLWGy7g7UMlQ0WDbP4sSXZ0/
aLcDKaAzRYy0CzSaEgILElEKRildU8ITElgmVlo2xCono2KhwzIL+m1k81IPuQONIXzwjQuQyXtP
dS+AVpDh+1lfZ2SopDMz6GQoPYTTGiFO/iK5qc5j00ypdWd0Er5OPgMr6lWNyzvEZFV6sdnT6ys9
RMp/nuS6EpVKWv4FZFttYMzFwaKEumDaqPURRe0KM9RzgYAkBH4SdQgyHKhPr7A3th5N7aM3IHwl
vpt6kKonaj6sUKV3OBL08SiQwQyOKvUj7gTLXDNBRKsIw6VQdR1cQ14QTkFzFD8FbnyL+je9EJzO
V248VVW2LArEbsHHcS7WoEDrGMAaZhuCiOL20Irv/yYxhotEa0iRpfqNeeYqfYgKr/mXVc2+3yXX
yV0pdC4Ml0L9g9q9HpVYPV0l/LrVPxPJ6fntjpaU7FmZhFMaLgcoPtIb3R6n9Y010bEGBU8ZjAfD
ixEZsMAz/ti0uqSYKYG9WkM+rKVyyRxUwkkWh+M/QRoteRUF0ZW2kohMT4Fmt2e5MlnSvCt1V3hS
kroypPDfCRaHNYlBntG8mRIhMLKmnMpftAvYs0wv+o2MsRcIasZydNUKn/zqpfv4OnSpZLyrVVKa
dJlT2xb2n3xGeMzsVSGiPxvbfyjeviHu86fjGDUuPC4bWRlJfu8Vd/KM+A9e6nigdIeSU1SbXJVk
gd4iR/4CXciBTJJ7byPMgFRO7WeUVl3lP3cbk3Zj4BMshY69LoauTRsDRi/DT6ay9n1CMwnKbK97
62wvFfQ4J1k/CJqm86Js1373lLFm6vjtFNajL1wndDTMVUjeuVEKUcIARBaHAgXp03636i7uShop
wWwtTaOIhida59lkc7whpuNy6kfIRunvo7+M5wd9Y6hVdyUoT7L+DAgQQKhpeb5D7kgdPKAqQqCy
2vNpG54wfaeE6BIjzEonRBd8OGsqJ7GuL90Zl0FkXhcU8vzK5HuJOxV/SeTZzpbjTaeBSVDUxnRx
dfMxxvDsFG06OGBI8NeMcn552UziwQxFw/kbWxqRNnK3IjKLhrNYFrOiqy31ZRF7C8Rd3zbyWQxW
is4scocMhZ15LM3K6acNRAxyMRG9g2myuzy0dNrShTTFXDRG/qdUboiplxLbwjro9jdxj6jvact6
9B/9s+dFEHOlyCwo+OFSonfCp2Oj8z0smF6hl6o8fma1r3QX6l6B5BzYz8cu7qzEcb/mao8VUKue
wVKUcLbbosTm2EzkDhGl7uaNNUvKXzF2XRkKoD4k1jwc8ZxdVZGGGWnoTQEc7VzibC/K0kabRm08
9t8Pgw8pq71P9ghDU6Zjl2DoIwLofqm1lIP7BBjzz014vlRFR1unxAz7Kg4XjpAK6ejiviETaiU6
1gTkNt4yUAb72b0TXtngY2ml/3/nok7LNL3lIxWuOB16FXL1v+BFuYO6hEy3ugFM/DRKmrwRP9tL
Nuq3TpWaX8ElFjpM1gmzjGWJLecjPhzLmKYef74QlZySmeCqY8UAeydMYcBoSuIkx19B2pWyolHG
zBtG52JDfy6wMbAe09aUt/vHv85EN2+cycRbzTIYXkuNft4nYFefHn6srr6BIX0tkP95JlKdWMfd
H6aTXdZ5e4L50Qv0YSnzHsPugzdgWLD2K9FVn82DHzcgdTDJDbHYwoSBbaKlzNEBcgsc0lWJfLoj
XD1cs/tL53ityYkdanrZIThOqg5I7/wM6tfb8rdlx4j9YAwRiVixUos4liTid0BZnLfaWLiRTDTS
//MtEQQeAhpVUcpio7sw5qoKB0/xT85yQ2ymu+p6Ova8RMgvrcM3Da+KvR2goAHLUcg2YLqxUhm5
3gWipbRAFyFJjy2ZoM7E9j8SIBwbLT8k5cthYEWCoELW9+rZmY5roF906tlWet+f3kCP1SK9M/rM
vY8gi3uYSvqrk81+4cy0Y5BnKxvbSuirKYGgazq7Sk2NYgjus8HEgTRbYv8xfZbnKYdmS4xHhvhd
ohOQoPpySVTAJOXKOEUQZJdtuyOQsxIU0UJwbWLzV93jFIqG2HvLoHNug5sADeOOBctmGBW04s89
NfxXI4K63UuT3K6p6Obw4EjX+DIOdOacJhOuECKhkoymZFATLTcWW4+P+NtxcWh11sIAo3+ZCgtZ
uonF0xAcFUYZ6s456VOscZ9Fk32sEkWDrOqUvRiN1WJs2UZOlM7Fq3BTaokgIIssCsPuyhVzprtL
sPsrDDBV/i6y/d8C7rG54kVFQZew7/1eGyLKpBaRIN9Rkrv1EtTzihT0RDJX6szq3vFcyy/mjRuI
XTfL8ZEoOBEVfZXBhnLPSQj9KTL2/vCqb98NjC7oKJ7+8mw/viqhwT8ayhd7+cQMTkveArsBKqwQ
Mc9MT+4Xrb0pbfgA7nJlg4a2BB2U24Ir3diMljGZ6potQV3onIK4taHYiu6rklvmqriMudspwdff
nYaEKIy1Hi5eQG8XKF8440JSMwmcMxhp5Pwdl1hhcYvxe9/Q8PCiqQOKME252JMWXtnxYVo3LZDw
pQEmPlC7aamoLbH2ztKvkAulQCZ6e+NjNuayS8AD6XWnhPnttkXlKq9LDAyZV/Elia3iTTRr24s5
QNuszlS+k6LseqsLBvX6Xv9c5Jb8wmqdBw06nwpEO0soaOQFr8JPMfmVlA0mmcl7vYf0u0IcCuDe
MCdk0wF0WFCm18J4hoGEprp1icboawOg6GALNcyXr661rdoUDJv/fz3NfBGQugYyNjcQJJho2ozm
1VKnRKADEXlHah09q4wdZVht0DHGHCiR3MuZmtGm4kujJMLpDsNSpi+VaJi8hNTEUEknV5KFm3bA
hAiZa8jtReOwzMz4AcJULwu7sC2+Xq/j8v2uhxyYiJwKWEYFmzo3znmjl2bJLFnS6Pgn+heRtFc/
AzECC8mC9ZaFBp6FE7bW9lCl4KUmiQTyU3fEgRZs1Hxcn6lgibNoTVrRDdPsiOnuiOJ9LYNWhwn7
LvfG8aHy1wRIPt9V1psCoHa5v74kmGdZ6QNtnpHcCswGlEC7ZpSX56+iG/qiuLtbHs46Hed4cddS
+LMfkhNrNg7obyqB6WXeBJoQORb8Vvrs4NfYE+VJdIONcn/iB1ctIpTmt0QSJ76gu3EB3j2jiEaq
WNpg0W7Gdsjuj/xv7RdEGczPUJwGZZzXBSivNLqSlHG2Zs9ctRmk4VsjUTOTeidlWy1WYpHSbznv
BJPOYMndvSy179IyVjW3p4TihdtdD8M6ELki9sLAzZzDduwlvtAEI85PTbS2gJ9Idouv0PXy4dap
rW5plxoh0piS6chfKgU64yGyi5iAmDpPkA0qvRbYD/ffokaZ4E22rUcrb5ZLveU0pW10StF5NED+
myz4p3KERuJxJ1ZLOgdhuOwb+pnYafTgSAyQJW/SxvUAg/N/F5vBdI782AoWMU1JZli08CUZknHT
ZLmAlLbD9WffI2GHXgKjcK9FfEAyWnAhq4vp8F5O8J1jKPJyKvsH/1yInlH0cLejPwD0p3tPjONM
7WcWWq6P3Wk1xLHVsCExqInsLxjvRo/AqWtps8t7f/IR/XTTJoRIgmzoOSZW2fg3452U6j48UGzn
gRmH7uWu9MzCTDDiL5SWBrXKY5DvNH2r3F9XVHe85Es8oXLdHtzKlVd9VWYbLuMjgjMjzxvwiOJf
qV34DtTTe+EJTwPwPI8fIroen4avhaynJTswqnHPIgD38eaTbDriTdM3jrKSEVawcrYZ1pRStOkl
Rkuhu4vtRM7LklIFQJ/DjiRXQ8LmwKuozfKKwEcwmgV/K/W8XXnE/ONTMtIOYKOzCBdP3HhAWgKy
6IONhu/njBjZF7eUSSpdsJBpdQcTuZwYytL2JYuRPZPn6/B68U62qaBLlykbufA3lPkYai4TrmSA
psa3e5PruwzaI3ub93+uz1ZG683ny+eiMSzgAnkCmuFlhTEBnRr3sRUOl4fhJhga53oxhMjow8uO
HO71YVw8AxJWXRfqYiHhTppWWtgME3dJaIwFiwAZgKBiCgkKfW4300x0Y7ybV8irqTD5/jlruO5z
5w/Xt8BqhbH/FNxZiUNWxZkpPCgLMGyhkSr1BfECNC52zk3zhn5nFC14TNALruAB2lqL0QWnVyGz
cWuq80SEGX+8/PhrIPl7ySbNl2zcogpezWB31P8nE4sF2EefN47DV+/pEisQK4EFYN25XJnyacMp
4dlOGnV18gteaUcXEDW5KfMTs5g+tM2v3ZE1WGBbRnboRI6/bnAxSBY95tPJJFxuruk/BU6u2Vzd
KDSrCiplWUevzrp2KEWWIhrVwXlvwSfKGS5hJcP98plNZBXQrnJcARSfFmevgya/50YGGXlWtlA/
XX17UZViQcgL88EQQ6he1orLHAnlhJCifRo1yVikXGPHx5MOE3dcBILFOP8EBSbc7lw2ezdTdsbB
aTFkA3eCMMkomEet6Rm2Ymr6kObUeH54WR3k5GqqhvZSctCqmYV+BdzjklGOW/OKhlBPEVoynPvs
zELA4Kxc4kxU3AQQyCPP6O8IqC214X+IRZ7kIxvorQFXlEDSEMQ8cP+ALzqu4TR8+dGHFa3Rq2rx
n36mNar+rBf6COMxm0NY7rdRbEHqtA8ER1mlnoD1gXHiq8dv/PENiRNUmoKuNbbAeMAWUUU1F4vl
Z1JEP6frYf92VnaUpTJeJOU2eH5uqnxA8HP2z6Fv90aJ1sn+86k5n+gOyKlf0xcaS+QVaz4jRr7Z
aGFbcyfbqMzg4QwQ/rZ7atJ9zS9jh5VDY57QdqKLd3SgNYCt0Q8PHHh3sDHgyfEijqxfPaJg4l7C
lN+47dt2u3H0DTuhq9LZatZ1dGx60IFC+u0xlc0lssC+f7X5sjzeBnFch7wHywdXJZjAOcBGm6xG
C0JiG8BLJ8OHYC3nLz9fe0qk0VbxtR5QxqCDyOwJmEQpjmS7rA2dtL4i8/i3BsTLoXTPr3G7iygO
YG2gH48gvLzWhOR1nQp+wE1Zt3/xH+xK7CTZ/CSaQPyk+aLbmvn+qdzzyBoOmAfAZYckwk0b8dzG
NCPQf6c6wzWIYFbszMuGZkq6M3hlnSL79rK6W8a1dkBXz6xxhK2+/elq+2Bd6goR2WSyimRvXLPD
BmmDOulEkZjWxuj+sbg7+TG+GsHici4zWctFhjbYNDrC/2Qnw+tB3QGhha+P8Zc0DmvAga14q2uH
d3FnZ1cRkOuxTyZhFU2bVpGOZxYx7vAbIqMMZOy0Jv3F7U4UHuL3WetSNkdD2V3bRZckmCqStFvI
+DkQpIKoAqSi45nAH+3Fa3sYLKvPttFiVGpC8uHTdDihb5wni9pDYfN/c/PvRuU1Hdz0UcBexptn
a8a4HmPMk1GeiF291h9TYsCMk9Hy+i7S7poDUJy5EQDIeRBP0FdmvIdviZqkxAiT1vtQLzIcL68e
veL5lxIM9iG5PbUzM8XrLvRgpO/5y/c0B88PW+0I/+pmz8uxztXi1PAbb7YCRJE/j2Bd3zw3YsvU
WTCOBzgDMUWYnCZQBHFid4um7zjRZlXHfaEQ5QVXqPDqqdKXSXyvkh3FHnJwLHlTBYmSir4OuIDU
cP/ZijozRdp7bcujlyOmki2rGjBcLdvNZr1D2VC+BGowvzJ3ULdRoNbIZDwJS/IQy3xqf4AFf2gd
gbzY9TbK4Fa0cyYUe3G6fWHDze9VDR41wTTbNLjTTcFwqlNl0IIxsXbvU8GHYPwStDkK4LAQgpiK
H8nfc81UkutBas3oWX7fz8D4EdFDoSHP2Fd4i2XkixnvzsRd9anp/rh/fVRBxzOYmXxYvbqyrKX5
rlUzQvV8wgSWkTmLvXbs3rSGNJM049DY2GRgubuKrLzj7aU/nW/V1hNEY7nUoClq/RsdJvVYAm2n
wcELtaEPapK2PjqsbbdZ0Jmz7/h+apaIrzntbBAqtPZFBXgzmkkOY6CEFFis0+L2bPmw9dmBiWwT
Emfe1EatCxIHYlJ8ugwIO4RWbYtJew6PffqJ4nNwAzyW9hgIh4mso8aubP2MU6rg8sAefgnnt08/
1LAFnUgvkKzITVgGnaknhTMuwk1BEV/AQkeKgAPFA94dK+LaCMLaM9KfuZj8T2OqwbEIF8/zf53H
XcIK5lqEzFsmtexqS5Sd9BtskzuFGFYmYjyHvI7QuTpmJOEJGllOZgoO5mb6Jq+lnK82N3FiC+98
q14uRr5FuOFcelUofKbd5dt0VFCPwKkCPxkQpv6jNPjtki06982OQMAsd2bI+q9PL3I0Df8fdAe6
vmNPl6GYs//LKylWN+j8Ci5twdZsaP8Qlcsi6Z0uYdaUVUxBhDSV4C5r5rcIQlqLKt+68N2JqpRF
l/A0vQz2hHYf5sitgd94+FmR5Dn7gR/+oPm4894E/Gnq46Lm2GagSUL1sDPl70aLvAZpSAJmh+s9
uLtgserKEBKqH/HuZ8NhBmY9Uu/LO0+KhgUq2DPmjpqQhuhnQTTdULkfBmcMHu6iUUj26xO+WSd+
6SCKBSK2hgGjcEzKby4JUEzyacWx6LpoUQsWKU2NB+AgAHn5mgOiLzohdlbegy0rnFzzmOxkrcy4
CQZQpksF6y9RP7HsU6yrSsUTz8I0lbIZXwOY4P2mRbY9YfHPtzn81mHolUXYsRpcIXdH1jCbttGo
Z43AAapZ6Em7Pnbfk9n5F1uf7z260LO1GJWrVnvpOAa3khq2uDyqQnzNPecb3trtp4+u4FotNtg4
+zwaJ+aNXDIbe/kqOKOPno31bSRaXhvcGyLAUYmPbUVbp28BLrOK9lW0nWdE6T1N97YUBm5ravLa
a+/bzv/+rTSbZrM0fhPQ+qXoch9NZ38MLH/DXTXmhq2SquAlFAKVcXPjkiNs8bbnyR7zVH+nhCLA
iIIeYPHwTW/h2VnhN0lb5/Ak1M8HSRhs3mIhWzE5hiSgxnpfr4FL3GbXQ9TZp79NrekZNYwm8X8G
TZZHBRXdMKOw5puXRgC5C0hBpWlRNB/rXOu04G08ExocGsPLCPDAGNOKU8EmP1jYlFL/OftpmJrj
QjbWLYO1CyjGUeKUJ4xpeT7nG/TkLCGiSL8cNaaUrcN1q25rcVluQ4RNyzyZ4Bo9geqGsY13Ne47
LCpjEQril+IVNeTbJJVj8IJC3jLD6ImXNE9qioITyExrLl+oQU0QX16DfNS7rphjxeTvHhiUqBtT
AQ3VKa/HrmTAYcfnHftCSB3XwxLwYrU+ruY+7oqOp6hUCx2I0U+iF4IBb6fZOouWr6IYAcT6+zLR
ABA6nwSNXzfnRv02xiqPdItivlr3IeogzwWbeQ6qp9PoWO9r57X+WRVxqEFs2MiZl3TVl/oNMafu
32LT9pKIx1E+uwKV0A/lUuKyfMsNzRFOhNwuTmTs2aSWbJjz/2oAoyJBGCOXEjlVF854Ue2cl0r1
qm7/PkaI3QYKYjkD4uxNJjrwUK4X6her0mQwIdibf625LyRGgbCT15GuwDyOp5iQpkW40bcf1o9T
B8OwXcrKSZjVAm5rrecT6kr9xa+hghxqO+hc/MeB4l9Qqrs08hWyQeZMSkjK1JwZow9f2O97J4j2
HUam5BGRe6XjzsvypvmG1hRkShVcogaitsGbM8HQqiBCU1goJM6xzRMBQeoMLJmiEtOxLZG7KjXF
Iq+7cTdSPzhba4Jcze85detLwTeENK6OT4miIFwcz61JWf2Be+q3/I0SEZa4PCXA0YPkvt3IyFwf
9jbNbFHW3VFNrdYDPJS07Fe325pAwwi5cEWBGJ1h3IMee5dT7f1X1VjUQsch/S4VXZ8nucijgoKZ
7KaiqKXOQp9uUcns/CqsPJKZTadDhz6O69vmvq1kIMy22jkuoFoc+UTkCCZ5GowVSXictKvUAo6C
sSNFbhrTuybgV+M0/ftniVgaJoSihX0ap5fXJtM2z0P0AgelULsMqErsxIILtlYERuIj+SNZ+aPs
ARYni4IjD4mUganE6ixQdlwFsCY+kyjTN5lu3qpN64e6mPvg9iUKGEUAhTvFVIa3gT0vHi1QlWom
8tZjK630LexoWTOqXDJ5hd5juTkSeMH0wgnn9JLzOSxF5Wwxh81qMVJOg4CNkvcixMfyA+3qfsgK
hP1QnZvLK3ojbLKeeOlhH7tPZIojDr2grZbsYKzxuQCazqWvN3frcDT5XSOzpyRrkGctDw+Bg8q+
mysC7USdcGdZiAZiY0L7ttYQ+KM6zZXvzOnEetadLl2oHoxVwemh45mvhNi2XAiKBsG3AWldZwdp
frlq249FfXR7kIQYrI/XTDXb8GxWodWkyRPp04qQi5VOruO0TMvn8dSAr+z2VsoVkY833zwKobTN
N3vfGXKYvEepWkMgs0YBeZ8BJFF+T0eKZsg9P4tzwDls646YnWcCLi6eiyNL99DFJ6h+ILdAJapm
apluBPzCjO3mh32bmVCwD1Rn3t4snrlNYPezKFxiLf53zs6HrQDJNLIUGIGf1J6G6aCNLPLkf5cT
4V4/nY4d9Gve7joTaZoBjKz47cZed4kkppLZECRK5VKxG+A8InxO13D35xF83M6u2MxTde6QiqtX
zBfFrnJP8m/m8vT+8ZoH4SLRGejJ7k+uiSBOhempTr7y0RcNVABe4mP+6tDY7pTG34R/Gh/C7S/I
ut277z2Eh7YdACfIrxXW0Skd9cnY0wNFJFu3bMniPLIHYDBQla/DbOL6uN4J3dety/zK74jJEbHs
yoxckbqhVtfD/Gupw9XYp/P0GMbNKpxIX/Cue/sevCvsK7RbdpyEfsmJ4pkpP4/VjAA3r6sl8Pmv
WMiWSXiVktDu/NEUHBOn0ffeOlbaqoCeAiiVEkqchG9bMyx1E/5j6qU46XgxmOHpFkJ/GR0SeP1i
oVo6HXBzdhggGxCz9JJT0G5AFBKD0CkRRMGcPEDzMiC8nI3cZdHNUtuszsuNJOGxTBZReqH5Ra1M
NoN8p+B5gnVZ/9ezJfnxwDjHQ6QaOQQ6rm02oj80EuakibyLQoVsejKoJ8NtNCKDEO7nQtLvuCiI
yNoR2kipRYkv9Ub2rpPURNTQdPDhQYz4C4ir2K5LYjZ1NfuoKFaJvakYYoKrt9l8xk7Jkrz5YP5O
iHZRm3URt3lshZXLWEXYeB2ccrSUDbYUri8IyoPUkiKWqGPiAm+IRCWrcOIQ1W1r226DXRSDHz/O
2KlWCkNZG1GodvNqu1GMe30KgYq7kaHF9uoIMjsnC8UYUpeJKIoCi/E+pGyyV3gciLpKLyBFXUUR
cvONOh9IsbfNCXpgqUUWMC8YUBbSxVfRvMfjjvHg+lv6U4DD9Kqw84p+8yJKw+bhu8CyY0dHGsvQ
4oW0g8RXAoXK0VyyReaTYbA0jM+n32589T0mUiN03ofG4CzR3W/qtxfDkZ5WoqIFlLZZt3NkSLDi
Ie+T6iKz75/cLRSVkx1/LLyDsrgXsuQsUqZBr7wOh3Nl8zn35ownZGkPE3/8Po4KplDEDGyb+mNZ
B0WPDsXBYtaaNv1cTMj+Zcn+iwbf0UI6pbld6tNdFh2NSRCMdPfhGRiFShpGyj1SRiVzzL9CVJxi
zhc7OhxVXXA15sXx1hvW5lpuYeB+Hh8SQ6cFZ1ajm/Q6RUefdnlUCX9SycThQIZSGsbU8j5cZ8p0
q7iDokfTvh6ADHN8VgHwh52B3vgmJz7R4Mo9aIcTzpdWkpiVP9xRZepg6lLPC+lxgLeCm/1d3nI+
iv3Akj6jj/atRQDgtvvBQTYG+C9ZMnz6mCtVCXSL5yGNWSF+5+dn0sypE8t9PQIsT6p6oFoMpr+U
b+ejYidCNBkmDo6R0cKvU4eRhGHljzwMriqJNXgf6RU/hVg6+NCAiYH8ELImOTEL5HooN96bpF7y
6ZtzE3r6Xqp2EuzDn6GlBcBPLqcdgzzKVUi2Dhe+2GwV1RcE6CeVh2By0/o8QC6TQFW0ppOUPUgd
PgaSGnXr+nQS1I74sfCRmOc/rwN4eoyLzBMS8MhXkjeQ+fN2W2/KDYkszS4TxAm+Mc5sVRz1jsGo
ys47qq6nwYZktXjw11G+pmrraijiLZ+hOogyPy5L2yyYkuk44ebR9n8d7Le8LGwZvznUiQDlIfw2
qaJuIDTLW28SI8c8bmsd6vZ9BxcLDjCUWUl+F7EiS3zECxT9KeGWMelgOwOjZZl6XHJS8dMe0Sq5
Nl268KM7E4WfasrvwO9EY3OFiCNV3tsfkyQr5AwhUM8a5kkcRIzBNAeSZZkP75606qvbo715qsxN
9LCH+77Cf+LRIdKJRoTtLFc/T46BAnoykNKgBMEby60IUB+RguhKe4orcaLlwgOGSl2XO5/X9pUR
rKKMFZ1O/WHThcABGfqW0XJZW5peZfZ9562rEfHQF29H6m1+iB6Yt9G8EYa788p97JP+cn2xtAyu
h4CPksXpgDDMsbrtsjtCnNqfyI4smPkTzM8y6IfsgiIvmJFXaEwtN1CLpuRGaw/rgtG5l1RS2u1q
16EJKVkPVn6Qlb2Xy7Eum6WYvrOUhRc4YNE4kRbKw8Xp1k/MnZwAePjOiUHd53XFCaETPxqQOH/+
HDFIX8vKfzlu+jsK7JssRSSsZ8oVOqTGS8HRtPmBdmjglUAHZPXTCsMXwLmwZCxWtakOgHBuvaQB
l0S/FKSXEcdex6ze1MXt7WlKaioso7TuUgEoV369Fa1mmuyo2ILdjM9WHe5YCS4QIM7gJRPgZqnV
1B+lmEmsMCFmbAcU4X+Gw1PDKkkqqPRWLy6xHUFDPMbGmNsZOQO59Pg7sYxBhPNbO7LgeWj2mVXP
c6dTKiaC5mitiGkFCQ5mL3IiOtpkdDJ5viB/eG0Gd6E3ISHoxO8jStZOPBOiIG+qMS0aN3ERGZmH
AK3q+QF4zWZMyUvbEyV8wnHwM+oz6gLhogZSVxOlXVaier53sbpibKwE/ZeBvgnYxxjLmx5XeCKa
oTmCHcLy9n0mGi6BTuvYNhF6kAPNE5LmEAbwg0FbFzCxt7aJ9MHg0IGYHlaRmQXMuGX16OQNhvqi
1Q/Up4m4y/eMemUWX7AJ2e7QYrN3LixwDxrGSc9lXqAp/ufVDJoL3JoN0C7vWVQ3sSLoGZDelJA+
AGMuRgifxPL0PMJIb+CELyqsdMY5Rt6st4m6zmJKLrBCF1rb6e7KUcHpcF2PxeO/yCEnTj3MgfNy
c+oS/9dgHBjYcs3OfPvm7SO/FwfAV1PGMNVWuVvC+7+gxgmrTbbs4KtGhzi4BV456Mmj6R6GWN0l
9iwaPU8QIGn/EmMSxlKSrob5hAfwmu6pYiGx1YhPJVIwiALSUUqzbEzeTb8zt4UiMt17RvEnEdRa
g/tBJG5vn1O7UiOhU/UvoP0ZtEh6kX0JMwJyqLmHVttyi95CB4Lb3oPNZuPKpMQ3EZrxSbt0Euao
nkCYFolQg+NEWkW4Q14sgKwAgnKZ3gdxTTnaentaT0KLhl/Zwb+a/YDyYNqMyop3mhRqa8IVFFnE
kam2qxBzb6SR45qKTH6lM3QqSWP38xnvxdMZ81r4OWDQ2ZA61ndEd729HqaqbpgE/dOnYCjatmTQ
I9qYe8ssBorEsgn2xVEMaeXin2sITBxPoZlRrPRVzsm8ptwnAyA5Hxs8CuvzspgYaOBOzC84SUpk
M8LvZCR6QayrY/nErafzwnpAq3nQF4RiS8YN1r2X+2vGBdSMme7icwQ1hEtDKWsp++xQ4Vl39Qrx
ro81RBflKVgAppnHy2BbYZJmq/gGDW4ttq4O7jrfX3DYZjJIZBr+BYDxu+Tsc61WWUjwEHQ+Hi6e
bk9d3GD/iWm8AU67KCYalR3aaRT0zXJJ8URDGQXmCKyR3w2lybrYRuOUlLA6axYZJa1D29DRlDfs
E4c+EpbCy4QsaY0WhfJLkF+QQmf64qcVcqdpp8jbbEESkerX8QQ5e+FEU0OcexkHTjVWFJUA7zMD
BfnDnRmVkKz4Vaye8KELYii4yvGuNekGilbEQ+ACh81rI7e0443Wu5DNMN14hgpG18JzE0E7tIrc
o1k5MQo/QnYxSj9L5uAXoxwdCHBkifhrWjUErn4lpp+VG+Rj33fydQ99ySSwB5Fs+WLbiSofRJ52
11CyqhF6HqoEMv4I69VdzIQrGkrs6GOw8Bnjj4sY9ohHcfhYhEVfrgV+5md7k8f4DOHawFDb8jep
1AevcVjQmlEp9RX/CoD3Taz5SRaumTJQ3XzX8nvO5x0N7G6fG2Y3OI4ZmNOoGVHDf+xlQgYsVx2Y
pTOrC2xg9t2/pD4ZA5TpZPAlJm8Ba6/yel+ILjTOeLeaf00r6dZHInv5BS7C/P6aCbv41nghV5VZ
r1HOcTJqIosDtaHn4lePtHPe8rAhynyD/pj3i8K3hBQqHEW/7u0vm4Omlu+lJ3pGKU1NU9NMBPTu
eZSCH5UderEkZDwLftD3u6bplZ1Na3Hrl9XxPiwcb5ccU07ywtYNE782iwU6rVzj0VSo4yt3gYNV
2uSMBA9sbEorRbHgppqrrZ/R+EDby2EriS2LLvnEH1RNzAvpwk3FzxUabSh/ILM1otB+xBHxsbMC
moNGN4uA87RYzf48EIEWBdTYdRrYpmlpeK7+7eJJW4IaECSxg6K1WEyxCYs0ed4qbkrBGBaqkzBn
Dy/+nMBZXmBVbbRWcwSuTFBQ41cNhNPnrL8+59hLMrVT/L1xwgn/t7MDSerORTXKls8cNZQp5RF1
FifHEZ1jra0FfJ+YIwjyPyejWYyFXaL5Jh32qM7u83E+BR0MdsT5v52fQF2k6wXTxE1jVRldrJz3
La10zxw505KydimEzYB2NQCH9btYBHhN0kWB8VFiKQihtoDy+p1AYycIIahPu+HmOtT7ivcjr3/R
uuiG3yYvJd8ucbqY2Hse8krt7FzdjrEPg7XtMdPo49RyJpRz6UooBRf0Yf+DRUJnX2QTd9/Qi3AE
tnRayeQZ4bQjCzmNYkUgbzrC/NNFRqUJ2Nrg9GSjltfLCmmHldtzNSVOgIX4Pgz2dzC70nXE7ggD
v36acoBoDtcP/ReYyqGRxE3VMcltRDSLoBZWuYR3CkGrhosexzACnivDu7jPNwGn0dnImBdLVA6Q
ls5vC2lDpEHJ8lzCacGMSoL5l8qyR5I76Ri6hErV5jpZeKGvKodCuaJguzFw6cvn5rCfDLJOmUQY
4GGkIJ2JRsgLRcl9x4iqiiNPLPw1Rr+vD9ZmVKa6C9w81O/J4ABHsc+Jf91mKYUnVKZUnUjj4Flr
oPc9sXrRXEsqhJ2T9YWPuEcTcKQshQtCFlv+ZaibsTJz/lDeFuU3clEnooI0HZcNYBT8XlQAOtqh
BpmW38QQgcUPkoh7SuXshOddVhoLylCHkrXbP1uDJ6GmBuF2eFcafxlh+dqVUZKVJHvnCS9kxpXO
FQgTCm7BwyJTGxxmMft/3pVQoWW79g9GkEBbgX+3WuDXbM5nqmj3mlKkVyqzl9VEAWiKCEArfZPt
XD+79kvszf7IB9e8P0viGq/3HgXjkWMBmPQ0ZIPR/x6mP94Cixfx3wxs6bRcxhqSfFnS7opqb+zv
RdkBsackR599GVikFtn7ogOFXJXzHPAOtovvqi6eu+I+LbbmQfwFZ1Kvk9OLxB8wPcj78fkvKp7U
JRC6LjHTxWo5KxWU1LkXYJwJbK7IzL9H0mgN0Rchx8eMgWtYyC/X3P5LrSHZzL9TyJo0hD/b7xWw
7i2E8pNYrMHSEBFpEI3dbFTSgfgpTncghusDEPYhN97igfiU0oApBAnPqal3EKae4yetlo3LpgjX
MbIRA3M8jCOOob9T5CmNlq4gZDjSkhc3xSdcuYgTclX81cjHnTculdDc7EpGiBihdkTVHmaf2qAC
SXJXcMCLPxDCN1t3v4ZTXwKVvlnTd9mmTSDh+gDHZa+SIumiDqg3CEqr8QnOLBIXt1TlAhGtWP/s
f4FM895BVZo14kkilLU/UrmUG6+perO058O+aYXTgRsA4kHGm5BbN5cCEiXrbsDFLhWin3cBmAhr
LHiGxB0/Pr9QSP2pt8Z3rcrrywmX4UJOIumqHgRMJKQGlcFJMS1OwOKcPi+07kl2H3UnAgyUCjO1
CXNl1bCNw5L6E8W2hSUwaEmj/rA6fl2C4/vYV8+qU2x8ntMQZT5MVgV0UQA2yzRqo2EMZyLsJRRP
ISKD/QLngjsfETy/CpWmR7yhtiBaEt2gVgCpEyRLOKARmteW7B32GYh22Tvvdz9tELAHBTMhqeo7
vjD3gIx8NP4nI4Fk2DNXa8VG1sBwjF5ySmzeC6EQVjOM+A34ZrNbxPffJfdYNyYniFWcBhx5DbZO
gtrBZlm+qAoyCM4euNyNnC7b3f3hLC978hG9hxVPFZm5y2OGv+wg3iaXILbsVwri0uQeBjf2CdBl
SBVe6sfq2xkN5zcEArXkK8FL/PVyrl+hOT3lu9EjZHVcKt0zOEkQ5ITPSjgrKy1IIvbJupTU29IF
3emfhc3KVy+mKIZS4VX0LVfULuUV/pjAQPrKpBTAdTwIImen+bGREdWcofNQHVkkigNT596yxOtX
TzynJ7GbNtvM/volhbBnNWQy+bHl4MyrDBi1uPQjIx3qaqB25wz/rdtdVHMQJlVdt0VZsLVcLd01
+KXi33jfMKJwN3A9B+K8ViTH3Wsr9W5PegBPMwPI6CFKg6QJ9HddW1zqijflXpf89VP0eJBu0yAx
KtSkdjmNLSvQXvdgqG6pbn4/1r0rJsnqMBtnTUaLbW//+2crf2gALuAIA97o8KN6mIGC/TGWFXPx
PXIkq+uk2isWP0UhNxvUX9eHSmfEZfw5V5rxohtc84+Ylc9BQL9leE/9MICNe2GG89KMfbo/fwLD
hveAMSzedItv9AGpj0wnwR4DTJ13KAHFCZju4Hbpq7M7ys7t799dN/h+Z839umIYOQHckX5olu2a
9qHFvsyGOJoTvhlwAGunesYJCjqhXeD8ot7j1kuefBCC+2H6CV35ikrBxFVRdNNh0FxJcdlizIpT
EpR0NYoIRueWnMt9El5Pp67nedulI1G+lu8Ma9CyjmKvpMsu2s4RxFeM7d2gwny8ZB0nfW2POQ8n
fKaWfOC+JO3+hLpiRVHms71HODCPprqq92fOPbmuPLBLFPf99vyOpkc8fu0NmmdpbWTlvjM4IMtP
b2EQVsogHkuxf41NE2zoEH1IT7O9qGmvrkeVYmgEMFYMLr8Uaf3xH7MhDwBKUrSIAzzMpP6f70pf
pOVZtarqOOE5d9WNRMq5rDMQxyRwb0sNcb6wkVZolG9OgHmgkNMIERbiUkfRvPLLqjxSepk9SZZ2
UHPkrE5DSiI5wviZEWObmK5ilYJy71ecpFw11eg/kHObUC3k856hI9hE3ndG9CJ6TpFyjHrx0Hfx
2uGXKv09djWe+zppuFjohi1pWCOw3zI91+32UVrwtrqPZJJhMGQZf2neLvOeDFgeHUk6HbljD3S4
k8I7GuLnOixB0piuXwhT6ZDJy8dYNo2UGd5bbdQQrm/1IebUuEFX5Kh/DL1ClSN0jSVva96fnEXd
pjiDbANoVVf2uG+xT/72aakzyOWvIaIsgC1azP1FAaOROtx/QskKlRvVatrW3ew0CyCOYnCDF0C0
wKZYO/Vgrg5MAGMI7enlWEevRPWaE4v03EMGWjVz1l27lS8vnhWB5dLYqLIYA/INlidlRRZYgW8d
2pr/D/OLPMwSF163O6XGmeeoS0yrVULGFSQR6tdDhVqCg9oTuKpF5xQ9QjCf7jRClcQABbUHB3lr
BS5cqf4YaBAPUL+2CX2U1mvClpOUNh+so8/YQWnnhl4Ow3HXcO3NNENdYwZNURtFZuZvzlcRG8Sj
Uv6b5iQ1iE4YIb938U0rJsZDHyHhhTC3ViWAK6BNPpTeXmx6OfOb7GAEHUatXutINLKbxFmzaAwI
GkHUrMVfOqI2innmsgvMKCbNTaZMn7tRBeJQdvtoKzOE2PKfFrqRvMsJXiKyiKHrcUV6h69Zcoaa
cC+Y3fgHHy0ZtDEdKLiu/1psatsNLlu9Lo7aKjv0HvVamreS1pZHnB49EezlZFoAwKljwuebZGBG
NWeLbA+uEfOPrKjYsYbV16AVKQvaL/0JooNdQQ0kEyJtNTyB1hrOsoOhX7ifxqKEDLgIZ4DlFDmi
I3D0qYhznvMCgpLR8ZEGJgB5JYM9yU2G+BTKnIH2X3zHWqq/cU6WD/6o12zHXRJ1qjqMQlBpGh5t
Q9EkVEB5fxgkTlZoHz1TQZGcVEuRalEDDg/FJUNaQGcZfKaiL2215W6RlgrjjvYXplbCxFmlkRW9
B/K5XXsg3qzxxNCU6yCCfkeIhtuyPC2YHnWSfljEO9FKpWFZoO5geGY74BH+D3GEZqGQCnCZ33sQ
kguTInrb1BorvB0heUiAIPfC6ULFzuvzty97fWp6s0/HScsQ/P8KBhLq1ay1xwEcz5XIvV9hcHwC
I99c9A2UOfmSnkvYQHOhU12rN7VeOmLgrlOSCwKtAKgFnITXEzBLZzhLxqEfO9PLyoUHFhWB5LQ6
5XPMoGiq+u8JD7+xzFUqYhgDRPPnZ1HpwkefkIoxnTZnzz8A0VH1EmllD4GeqqQdWuHR0WgKPWFt
scUw1rTqH/1J2Oar9bvw7W3OUos8ktrBVfYLNS+goKD5ZH7aLk/1AHKmv9fJZK89uto3lAg64gAa
vNwNx1Xf7j4SHUIXQsBj66iWMe5BRJ0CYbBNO2J5E80ihE/584s/bVTZsJhi4urz0y07MKmf44Ai
mvt7Av4vilHQhkVSPt9TXrVYYf6pZ/nuKRbGai5xfx47ceB7xmHIA2QebiI4NB8Kvk9P1kvGegw2
UyaRYP4kcjBZlix3Itswj/ZlGTiWuZKLT1l8ln3VXPTlCIqgtqIJ6Ytk5jkByYbs2vyhdQTV5zh4
hPSljNZ0ANvvdaU/53v4rB7Z1aaaugktbQethUIUb02KnAZisJu/7ujzFO+HqJW3jSW6ZHArDFHN
UaMF68I0NuGdN9Fd5Ui/UoAG1TcbG9sFPZmKHOXatNuYzKZCly6FESSFpfQJHQIQG2hReKNCa/F1
QqC5ZxmIOjyW/hHLWynzYFyU8sX+WHKpldWEVLd+v9Y3WevNS1ZraTdAGUGvdCQPelpHe/50uic9
halQg6SMpfADWP6Kb66p1jHb3kbITkpm14JQf4nOKcrNcxQf9JSFcOcI7IUUiMulYkznxT1ZBRcm
QLdI1UlNbjOOFup59m5fsWbh271i0BZsBYelhXVr6FjCV6GHICihPKs6IDxnlm8jUsA7sJ0C6W/P
xlURJhZHZ6fDFdbQNPZZOCeg46Ylh5dSMir2QFGp3/LXwoVgcvoFKK/nApbXqtZaZcUZQc8M+stv
CODFE7ss7UJk974+X6xsmUCuFb5qMGU22RYGCkHYeWnlpXHRxG4OOt/exeJ+3pn1NhK/zUF3lwoF
mdLXVRd8T66ZIRpX+mf4JNrW7TEJT+nUV4pv8yG6Bun1PACmcT5/nr97B21A9eoUZhGEeohWftJK
9BZVvI+6lrw5okwlsI2+xNTShKX8o9N13vGomGxeC8lxmnnYlOhS38sy6KnCd8uWk0HAXYH1iYq4
SvnLBPqjp2TNkyP0r2RGMZLYxDyVNWpilEDpwGlbhHTi4LfnbgaoLRFUCUXG4rIPsOkgrMK4QSQx
zAO3WZT4vpTMVyQVTP5smB0RizuJJyqglV/AQOe7EuPifbLpzLJPb5FPNaXMwNWrckoWtHfT8Iq/
jDmrNoiXRt0r791Yd3SNTv3EQFHnq7/HycGYIl47u7naFLrbQpBbbfWoS0J55uv6E6IgjbC70vLz
6vFQzzjy8lyFNTMw3TW6LuRkmulRD2MwMyw5PfEfa8jX7UdKWrT1LBWATDzWGujD9LpV6eHWURLW
LNcxD7IxggKFV59j/MKd6Erg65O2dNqkB0Yn3x5zMo2jT+Xh1qVAKphxo8wPWHfSX6ECc2vsuJzY
ncnCOzMmxE2PpfkDFmgUFnoHqEkj5w6avGwizSnKWdqHQ41+OvzswZI27RohIHXg9Gg0HG3KujnE
5Ts05m0e8OEBMH/CxN04QhWBidodiKjrekj1QZz/2nfNvwJXvCP72FnyazxLZwow0Kjc8hvivYAA
Tr56khabPDZDKk/L335CAKQybdKFUBTXRGOHdSGyaD9UOn4V07bfDM+wWQQf9l9WNLXFMKa5jgeg
YtqTiUC9FtXsXWw+weKz9+5fFJEkNfmCFnlFAt0K7WC30AnqToSSst1mE718dRIqT51YXD0fRC8K
aXhX3cpkzIEoGdHp6cArKn8zfYytVQEmlzsm7VMofO5/UVnt1TmcEWidTEHsbVCqM7BD4TZkZSby
2c5L13PCjH0qe+3+t1bTAZc6RK5yLQuG+PCYV2L/mPThbYPUBEIs2YQWTGn/d+/NgwR9FLUYTdgv
UY4iRz23TbWnyMb8d8bxotsLd7EAaFT0faghkU76Lxwta9I9yLCAoBvOiUGPiJkk6CZzClUyRfe6
ff0H2+f9CWd6Fe1chHFIWj7oks0Oh0aBiFQS98pAH0On3KTGdNlLkv2B5z+Xl8knDUvYaF+K2BOJ
fMQCkBFMeGFD9+1cyOVcA2njSczrdFJEN2IMI4aa3K4AFm6MikZRI5OFNoX04s0MDF4cGSxImXKQ
lm+wJbRJFyLGi/3fPUyyWZeLithVegzTrIWq28SgWTqoH8lLC8z3IvWZp/OUsCYNUrcUg9DhpdKL
CtXZkhTlG6oupwLWyAC270hmnAxlMORRqSa2Of2dC3oKymfuyT61pK9aLC1VsKcLsR/gforxS5g/
8U8f8xpXFN+dyw4o9LJY1IXMWH33UQExQlaXmQIGuKcVH8YGffUHg3oSBoUREBIFxw56o3NuaTFU
GRS8QA5vlnNVHwMgBif4tUdDLosXL/N510kMvjTodWTkwb6Jt1XMTDHjcYvOw7qCpB/zDs3QEXuh
pYZTB5l9mZ5e/BJpJbqLmeo8gEImiV9Wull2bJUQP1v2tUn4wgB+l+XFw1i6mN4XZInj6Z+XKrbi
fZ68aQI5NEJMdcgF5hb5IOj00Y101pmwiXV0WMmSYvveig1Hv9qNZ+fWXQDpuM+QqmfLp+EIpIS5
I5rG6xDZfjNpGaNyj30SWKzWTK2v7bZJJ838ehdCn4I+/UVCdWlmVKFgGHJUyAOJ5Gy9J2b4hwtZ
e1lA9kpj8CAy2S0QKPV/qSVOYeGiwGcaaJUfraJQJNQC6hFrkS0jtZiCHdvCoqpPxYs69Zsjm1XP
m93i3PA71ypXkFKTplkpp8sRX7p3qQd+842d/SWpXY3Nhp3rrth4nXRcvglGx/lWr6C5QARV1qJ6
yLAlrwBRhpK9qVAxszLSBpahmg+rDrs5pySwQ8s0SIcRS5EKvl9w9RUVYEMjwokrLT10fll+n0gr
+tahNFtDNhqpVCdoJ6iT3TD7Vk1Rw7j+A77jaedvBeMnfRyD3VIiCLrqQtw2FB+civRuVU52VKtk
zZGyU3huF6UmDWjU5C6TksF7N4vyeFupG0IDqjNmMqXeFAoBfDN9imskhHywzo0Rc93keZjlGUcx
dtj7kyi9D99IJWtyUHduIe6XAkdtEA0Os+gvR7nj/cDKZFRD3ZobpwPh6yMIj224vuHqHAN8hxSN
sOcTPIRjiShdfe0jkHygYvhtYKq/+TCD89C8tqgTq8avqTS9ZXo+vzJDIojVWC3Rat7RLgW5GZB8
cyUv0OweEGArA7eO7enMKbXkUgyG9C5K6RftUnkMDQKAsytsb8zZcFyYiJqHXm3/9HXdcFkM4H7Q
pHHUtEez0KhFMnBLoiAE1+f9Hr2v04kDJsaDi14hjnOsc52EmTYy7scx3haaL66m9LZYYXdUfqsZ
iAuBNNg4d5/Ry1ijJZBcdMPp21+apBGmBWT7RfWI4TwOQL7SNxVXV7pv4YN0L5wGkal2gScfUXHp
/EuPQCtGyjsvJ62hgV4klmXuqXgKKJYqi2dEKD9nYM7vgTEdPhDqoT5xU4k93wPeigxQlywpWkHl
GafrnftRM9kfooyL7V8ZYv288wDwaxdXxcoNpj5OOnD+jSbLlsEmPZYYDH+D0gH3pWBeAWSO6XSY
JpeujEBUFSlU+0ycH30D5oTSMGgmJCyJf+3bzHIeDLDibja6ixgtt7mWw1vsXpEqfhUDichQ2saF
YdZyclTExjkuNkd91aZyXgk4DPcugq+IXLvXiW5ta1rpXkBMqmiQ061B4XUfv5MQE8TbawOMjtSL
saMW6jl4W/FDOTRnLsoX2kbgy1VQid14jvck/bQJHiqGurK7NRfeYBBHR/2iIA+8wTYC+62/PEWp
KkA/RUFTUXfh8XNcR7qwnseLaGPwcDtMuAJnQQ3WJONjyEO9KZhkanQWGAfSIltpQ6xMs1pMEBEQ
Abb5w/fA6q40Vb98ZGFXpkFeVhL22M8/xH6T/BlzKzl6AuWSRAV8qJbddaYkw9u7rwKdLVzIhTpJ
FkIfIIFHw8gKZn8rlDJTTuyfEodmjcWDsfUEspOAb82JMjSRvErb6rT+n+6ZDiXc6aTPT5GdkEVS
lZLfEcae8L/g/lpFimayFDQiIXwYFxv5vWGrui7+4twFBF+0we0rYFXSJSDgsGSe7KVUwjEixMHJ
1DGLe/1Vp/eRqYiW2vSdz7w1dP9K/w8hcr7/x6LtM2M4s+H3KDzwmfeNEMTZ7bwSNgbnLQ18WKv5
6I/laIFu0bcVauGUkE9zyihlS4yp3Xts8PalqlYbL6cJHbI+Lqh+MiB8yvCB1v7PmGzXLGsAu4CU
xF/tbrzA6AXIkYkLkpxi13Ca5cpLgX4u68bdVHZVY6YJolpfjPPxh4SnxOQ6jiN574rBK+JJQOpS
RIY2taFsPRfA1dc4TYyIiZgU6DCw5AKbvJOkezZlXpgnV9gYPnC2WDjjzDiTV/ECIJ3aOFHIPPq5
fPXrnsTg2TLutdrbJ4STcKnSvGZ1QOmiiDzpOZmfbujtKuunbiJ9PEKOknC0/KyrLE1CI8bONT1M
pHMNhH5fu17zF8HPCKWDrE7RWDxV+ipfLZJa6/nk/40OCJ8FMSk473M3X7ydsZNbl/Jp3UOu4VEL
sh8QYGV3BaA/uo5nkog7yHvUam651hoySPgFlyVkZtJt/U13DvWqZgFqqB0vdSY2JWB+IL7Syx49
Iqi/dmKJ/CCT0PUswcolf38QlI0nQGAIsQQD+mVZAKrr8It5CuPKiRtZuKzHImVQAMQYTlR9BP/J
AV0hlMoPMNmHMPqhtL+rJ0iXS++jMbdyeXlml4TLC+Lf9eVCTD3FS9Ph9HCJ9lB4iMQxR8sVrKvf
mtiH/TVIyG9qcbbzq7bNLogXJKUvzdBz/WB585gvadx+D9SGS2LL9ezX4OsvswoJDftGSMwS8/P9
jwJsU5CjTN/Khseq7unPMyeC1y9tGXhHV9TVHzcbFC+HqJ9RXj53UapzzBuBPMATeHmcviqLuoZF
dfzw6GsnJCKgm3njwJEpVp0+dbmE5aAvdSMkNUyVYmp+K4mZRQl5iFWZUQkkbB/Xt2MFyBCa2dpt
+6sSzaglZ3rzxQYWLaFqAIwnC+NrKjsob/0uKMzXBckL4CdWYlXlPiPhiO9eGodtYcmpyTw0VsuQ
TxQmYmq3SDfZcWPBjBeIjyWaq0jxDU1hY+u/Ybf+0OCxxIoKHv13AdrW9oiNsabAxfjhe4rls8bH
ZaXsyv3vjM2E9jyF3CQOFfQ6omumffmzJSYkD/+/989C3dWLatQlBOBGEMBoJ1H9cX5PKRugh3gr
sV/ZTSr1V1xs1VWin4KotznK5f1rhtAfKSmpNwWbOwpyEOT7tNLiL8SWFa3ZY00i4/ZQ3IFb64ry
ZlsD7d5hWjXDPYmOQQnPQS6AmSGKLjSSjJJx4NleLGN/HnlpzFfAmT4joLBxUxRQT+Rp0HJtbmP4
nXqns8cgw+i518izwoLuD/pYFYpnKYbOkBJ0dFrnD2bE/lM8AdvnmEqzhL+/5IrTwgA1g49aSeeq
lp3DQcZcIEpgcuwQjZtO3G2/QHMfr4UkM2v3mfCEd4JnjaLSOcW5l22XCIOVEe8NgQQfrKMHVn1k
5OWzUQQai8qJZlCG2a9/CRgDvQWhVoqYtexrFBYTvcvT7ojwVc0+UMNYCxi2S85+Eey2NC3JrKNR
lRYmmNCSBOfRdTHbRLxfSG0M8maVUFytRAn0rvOjK2s24Nizv6ixRgk8JGKaSImcmSmIb46Z/3XG
Q7/2e/YrKKY+4LY3CJEi7s0MJQ+rD8zoAm/2Zp7zQd5am/kfNmPZe6Qeb5RFNOTKgE/Tg/poqymg
QNZcrAiZonSeZcq2NLYvCwOaw0nAX7n/ySU8P7/5XJGGsx/DDJ0418QQ7jErQ7FgnkrWajtl7wd4
DQcYrjKGW0j0SLjgCmVgcXFZtEdhac+axFOD2b3POE8vaFhNMn2r6EbMu30J+6c7szpowlZe95Be
pf39dllTfjsQLV/ZN6gr55NvrIAl8PvDghGCj2oU1chddO4ql0xTT+WFnOhV1AbiqQ3AP9dpnoTR
KTemyNwINYdylsfo79K4GlStgaJndCwj83Y3gAQuASpMb1tXGBTwhbORWrfS7m2lgRbp9SCI1rjs
aikvknhRsnhnrDNfzHupR4Ha5TG7pzpwgnh7PR4HG2WIXblhIqK8MicqhCzJI9me9ucfnytRS0kz
NmBb4PZ7AC7n7Wgx6iZ16fZB2tCLTuOLPpw3y+vOTE8CCQQ6BO0oUWEGM6Gt2xQF5u3szs7We5B8
keT0X/49bhY0G74z+JykCHiE0ZS3PD3066ky33lmGV1YTpXzRryLXZfRk9Ez1OZDn70BUBruMC7u
DZXZ4ZdEqQZF7Fi8cWXg8PUNUMiihwW/H8eRdC2rnXiM/0bILtTiWCGAJjTUyNqXgYxlqP7J/kSj
k2rwgnFE62t6Ht0MyhQVlUUOJRBeIL3b6A/TZvHWiCU9jeYwmQrVNQfIr2m9l4IH0rPkU9OvQ7JG
pxgv18nMXmbz46ygpw0XyV0Oac/ihCkXrW0kvdVTfIWKad2NRxB8e7WL5qkGny5xMu7nYhKjKZ8i
lqANtz1UBrcCa6kxs9CpUjk+oOybkUcpqXhbRXE4B4T4oZRIbEY9TNSvnaIw0GG8IAk8riFNqpCV
/MMocAjDdbq6kkPZQSFohTNkg2jLaFX4WH+8k1zqotj3NBY/YSizvu67NF2tcvBlnSRBm2E9pf38
VRlqQB8UzZiBAjhspm5ewfJV55ccGw71AIqGeCcxjN0MuB39dCSN7Fcp1tv/Ve/MPANGajfVzUTm
dUR1+U6F9hSN+NfYzx6vitjjkpbxYD0XQ5WEwIX9yyyVVBBxB0qIR4321F/A9iKtcsFTpGxyuY7B
o0gLqL9yU12NmP5v1okKHhXG2f5UvQ2L1hhyuv0OwfQ/eIPv0B5B47u0Ml6mSQBCainPqrcRxclq
9yTAI061F9VKOdZT4egjFSkYQFafz9BkV940v3TV53tTTcAItq7lPNEtH00XIYqDgrmD4Cvq5axb
6J7vzY9S25BKCF1DFUmR794b3e4xq6bsaAj0DxvYBOpY/3CxUPx8cce8/HgOOMf5tbo1Qb02Rv/v
rWgwGeIIlq9sz9piGo8D1uZCC6RtLTH5lJSEzjG05/tQGR7RyotkvQTS0aIFlxGKyL90tuMt7oF8
VPnvKLFIuiPpWb5VcG6hU/pjjDJQYMZ9yUFlADT/ctHF9HYqSDrvW5F7nHUXFyjHJ4Mof9hYylAZ
FZnR55O8m1xOjngpxv0NceHMdZEUK5TRH6fh/XfDUCDTLf6s0UEEm4FYhTac6QcPXox7WhgnSGrd
dStIcxbkJuEHNUQc4xweDGHadgjV+e8NX8Qml6XNsbd1P0lDXKsd00qAFnA1nm0aTtI+2m2YKtS6
jNKebwfCzSJAxP5kVUMYnF8WEZ/aMA8tc57JqHpwE4X6VKvR04z+Jiy6Wz3KvFEWDmTzoKvXP8eL
tM/dQ96QbKliUev2YC9eVjt/fyFAdi0IGmYj8+pfu0GYSi/cvI1qA2ljIi1IN2N842AuCbdTVa53
qmGBUj6p9jJiDBmiXadhp84755FoJifsvgjAWR8GG4wr+mW6S7UFo5L/VjeDNtVZie8+UBGOBwxG
y6//xjJPkf+UFJsCA8QO45qqt0tI0UUpHyRBYnBOkHTjOg1y9W/xthjyUJRVIZHzVXidBmAsWYBQ
u9+uE2ETVtOBYsg80/H3AvE25axcN75V9qO0h80poYCQ373sFDSExc5ZcZFpQoUiFmFs1PFXJPU4
I0kum7xWn5euyoVU8nQBetXJgENIetRfBu9D3LArqw/aMjamGkGs8TR21po0bvXenbSLf5mdVlHC
+SEjXd7AuhVDAGnIXkZ+Oq6/Q7uaQV6ARMXJgUxY2evs31gH5VhFB9tNbtvK2l8RTF1FJ/VVzy8E
w3kHEcRKeFoVP+E4ZL54c1ZvDhro29ly1m+cq7TvtgaoNAACbKkQOrAnPYkTLCXVgMRCYsbqwZgc
ai7tdR/C26S1kgvJnRmRJk8xoJQHMsCrrIylIyosMTaOqOHy03bOG15lmU1AQDYu4AiGl6EshOu1
4RVVIuJUcnKx8XtTMudjRXVPU4w17oVrWfRSTeWJW68wXShqRWqINkld9PBrtzYo0XM3K+M19xVf
Bez/B5R+YU+Nx+UV53RIezo7VWwpumt9cDJ9Htqn8hUSUdjgWnXKPGUFR9DbIHodZhPQ59u27qXf
zeKfcI/OxScIycLFcaq3Jly5jWfIK80e3B85ySVx/cFt65BOmjoe6D48RSzXPkEWFO5lc6h2tybr
H+dkzU2WUKU1fxOdFMVPKbNWbCV80z9umsZYER88/eAyGgLIwLb80ZyTRVr3bsUXkO0abxYGzya9
FCWV+8Fzy9sOOqGwAPf9A2YVSxIOAEBT4BnJQ5qhSqa7BEtnFxXMKFny/J4c31T2ErmIqQAAdVai
mNDAIaEHK5szJXt10vu31m7M69uyo6thIjPtbhQXYbZ3Q4nB4/2mv5aY5AFZwy0zuMSltP0FnjrQ
salO8irPVGuzIvb2AG+X4jIO2ur5P17745BsLXUgbB0d/shkkSe0erMXStBllkpKGWCOXLldf7M3
XgSmugmJpDEWEmhDekUr43c5E0aQ37AtZV+YegGQJ6QTiJEI3cpW89lEU61tSSJ1qHo3sPRSZP9o
ELtVL7zjlHGeDjC4vE0B1OVXSD+MgRDeB2jXCyasmiT8JUoIOK9W4cqpLXF9CmMfsdvy0GVtT43c
r+7kM+R8NFUB0acCFrb3j1tu14V8ov34pNw/8odbuQddR6xpazRvfaflkFuvwesrbeUjjaV690Yp
nLJBbnD4SCrFis1e5e8ervU61/DpxCeo5DnR94TRjQuxNGOWsQPFnrorjM7FcMhXXprK4nv1CGeo
gMWuSYYeNM+HXiW81IwXJ5YWIsXgmJg1++NhXxp5gxouVEOXA00ZvDbbmzXXa6jB5am5CXBzrKK7
ROhvjwOwW5jRQ9i2MQFKGypbkOGZpXRfmVaBrN1OLkf/lAFpqd4G1+DrJKxPz7NIQDHw7FIpZjzT
pyImzB+sYQz8UugIknMmMIBz1Td2IVzL25VQ0GvX5JM9HRempFnYslTk16MQPqO925pk+Qo8EfIA
ADDoyolPYSGvOLM3HwvE1XcjQHjc8RsByZgRZlucPKFSSBbV/hytZutQuGe2HE9ilrU1sMKBETm8
dwQJGQ6pCMlM++NaPZliZOFLIEkn1fEE1R+4SCcyCHgSHTk5OhYzs3qkTmCyyx9mQZDW11HriOFW
Mdfb2bNc0A1h9A5O9gUNwNzZmJCCOU+OZG+ZrEpBVSQzUFdXkAYZlEFDiDjZgSF08gRsi/amU+TC
Co2idF1rhfV0bIZcnwG7fPh2HuK70qJ6vBVRmPs7bwvOifdayGQg6irr+H6Jez0jq1mEAPlsZ4YC
EH5z3NUmkgmZ9JNSggy1XgdGt3T9ACYilpr2dF2cHrRr5hn4Qc3aZ3nyrhcsiJuPyH/cZuHHdiPw
3ZEz4xxsDKiCUgLsPgYr2iBNMBSzCTGuruirsIVvk/bavREs15csSu1rojKclN0oS2JY0z5VTJti
YAjHNlZ3KGMx8Vl0TbkybdyuqOWXAPnZXlrnG3xlGxwgl6x8DhOVAhduJ3K6iqLGdrwPkRN5Hk1H
dl3KRYwuBv4Btt1VfSn+mNsmnho1N9JWMvkCWH82sWQQRoi6fwGQFryHhPGF+nTlZbreFnhHcPs/
YGH7bhSkz3H7esmuDHkdO20VCig/IJufiUoN/G6kgdkfZC87nJXyDnrMxSmfR0oJUaPy194mU470
IAc/xiwLdgnBQCCWgLLWQUDCgjNw8hXTUQznb8MC1UJRfmk0scAMnZPzvc2Zo+Inck3z/Zyy5agk
J9yu1OGVsePSf7EvlyUUuLd2BRa2WiNkCTF7tJwn0vX9CLIgeD3rQJ+teFPffilneTPdHUxO6zlA
AaGczpO8qNWPI5Eny2/Xmg3VWdVDtkMbaqaHfmBgsuUXBLdoP+opfbksJjaTdHed2IAjXeyStvCE
KFjryFQE4YaaY5vZqVyh8bZuqWpVoVclrMdMJVQuTogb3x9k0xFpOVsVfqMCMOHeasDghXl6wDYD
QNPpOXSCaoTfK37eHDUCuU2/RJXjd2yYpU09NWQVzITET5pM2sLXE+uim5dx4uCCrc5zXMS48Bst
Npt2SzTy3Ot5Swo8kJUyLfpveys7AGTWMuvIOeMHJsK2QticW7lNeUcNBAmx1reTeTySUcGjbmHw
1ce9wHwdETIwjMKpMIzPUSS8QaoPK/r8eu0XNiuUdMPxdueAKPDGtQ+XZndo0llb1yz7dUjvidre
jg8fp3PCxDeBIfG8aTZab8jFD5bScBL8w3FDJXG2QE1ys/ziHAlhrHB880Uw9DJTrujaB+Ok0T7w
uw1ZL0v25vyk5P9iVIsHIPIK3ZTKIVejAwGsVzZP4ndOVwSa5XSO8mi83LJAo2H6bVyGQvDYHWIf
JLtWrTZO+besBeGB4HGXta87YCR9IiaJZjpqODstspLP5YV2sioSLyDs5mJCrElY/2ffhYsPwZ9s
mNj3SY2vXrSsM7kKI51xJ59aXmWv5gcsvumrao53UDbj3K5zI+U2zhtCbPYLutWaW59t74lAC69o
GXWeAZh4UN2Wlif8vBmn1/xXfRoiF2s7y3dmJnC8Zz33hxhS1EdglmOMwrd8XxmrX7avs7FUl1mG
Io6Si7AogTt3mTIWXWdCR2ldg9C1HKrIKLecZNQbk8IJPTdDdRYsUMtMZqzIMK2vld7yyhFOC+hZ
RFwUyHh5XeIFfyH0purB+i2jbcvgLK7wOSkxlThmMYzTm7NOzod2T1edzTicnPLdgEoWbC1c3IdH
+9Numy7g2DkMdapFlMzXCozpVTzcVxHgkCOB7q4PkSmUGwErLOx7oRNIJ8fOcuVwVGrX4skeL792
wnuhodIF9cIE/JZYtqdg8QG3fwaNdGp3dmYsGF8mfrQuryD+1LuEUsmF3JrffO2Lb/U5LR3UBqtp
ikO/G6NIf9tam5Q54l19xwPsRNpF7chmEARdPZgzywm56MOq32KGw8jMtpZJj5Nxmj/8LYTw4vfI
om1qIrKIVCsNbhQlb9Zz+CWgCd5CZ6NXDnMtvnjbPAACNTuMrQz3PQQdBFgNmC+M71Eu+1SCxcJf
2Qu8bkxYq87iTNNW9FKUJeDqc87mb+hV1akuXelM7Fb9oFtAmze1lL2LPB+v8cLedhPaw6gJbDd9
R0TKNH5PQpVrSmNrOb8BDD3hoBHnC/fq40JJIAih20su+55Ocvav0izCuGQN6RzOcrbOqE5FVyRD
cNyCDupteEcrvS1pKneqcEtX8wJPKlPG0T0mG/cThl0Wl9NFvHSSG9sf8uiSeZ92yzyYpu+ZGflY
tuS4iN69vtEy9J4XRUfpfDqNdiWKa7nDSiytZsEP0geW0hhCXnZgzihZQwHtkza63seTfeYA4sWm
wo7GwXUQIQ/Ctiyr/jGDiJ8YbKaoNvgSUsufD7UEgnGPKKnMl4jTDygrrDvyb/Ug2zoUUTbHZiYH
bAVG7kVifZ+mxEkp576tR5KS3St2AW42XAVPx7Dd710cYW7aa1zeMKUuVhunDYHWoRML5EeYqsAF
xpQsr17LswYPW8XHvHkaB9wN+9TeYA368vLWjo8uQ9Oi0YznbC8kv+ypA0k1AcEqMEzLY+5IPzWh
cyaPX8ze9n6RuwgcmWJWIZk8eRyj3YBWGVXxUOyS3vlE5/JbSTJbcCRw0Hkb5XqHv06Oei6VlVks
pzKgUUjg0iYZj7azfR5QKdxEYKyNPyxHod4wAdzD0f2bicSmwTINgN7Gv+JSreBi9qa25WMB7Pgx
32JoZQIhbarh2CEMBizlGzd4bJDnDqMV20i6nz8VEzln2w617VnvQgZ0QrUGy553XOMCWNWyKZiE
t6gPXICtk6oA7WzsbhLa548PYb9ZWqpKVveF1dSx3t5xJF9kuQMfSjQ6c9SXVjZjcqcKbaP3sc7P
kWYis2XX5NMl0JUxRcDkcFrB0IHr6PX2Gj5CnExAB4AgBG85qDORjwrB7kPTq6Yz9M66BMRAizFC
kdS6w05HhlCIYE2xNakkHEZVV09qWnx/K0RNtZZ6EDQrJ1T2Yq10Sx4ItDFpeNUkb+Djw4W0mhTt
+r5qgFKuGCxrP8h7+CEt50dXuQTtfUCSvjEwNNNQjodDC83axSN4LxRWUYUioAw8nvbUzxNVSk+N
sXnzwRNPh54TBSluGSS8PoDO97bJ6XUL67Z96iA7FaUHMf+1klajOaCb+mJFNZxNrrAHitUyvm16
1wuD4ZO1tkt3NOaTXs5sqCKgrvhvvjB5NMkuyC9k1IKg45fAThKtWiLsGS9EqD4vt7XDG4w9ni9u
yvVrXW4T5uRHqWyP4xLa33D+sJSEy+Gx5sTdYCo5MC08p9SBHFoq1OhMSWJmdh5l1q2EHd0kTkJh
aAvL2Fb2ClD3aQ798uBN83m6xO644uLj2ycZnrYNI4MQHp450hS/NGmu9QcZEcyMmeiWvXVWMnbq
HJhMpvvT9mW0Z/zmwo8KI9wPymRYclW5v3eQEZow/esWDOZlo9p0tY0yHxMaq+TF8gUMsp9+DNcj
DXP9DKeUDX6aCA805BnGwsfFiXnUsY8GwRGWAmc6RVlYDdDkK+DKhA/zbXlpPoHMZJ4qMV5RfrKt
tgTD2BKFhSCqHuCiYwMHfqr1XIguRj+XFWfwbyNxDHEIuqzLIe8G4ZlYzQBo4sfsFr4noWv3qy5c
NBTesGPHEzxgwLQGd4oIE8E18PDcTzkchw0tMUORWiLkU7OU3Zz5kB+IQ4UocLv67kSxavHohJDy
nqJLamQONNN6rVpsFrJvFs/gX8Q4oUddEw5eHCLiY30J80ZLMoIg95r99+PBn5Wsr9GQUS9BJUED
Xz/hPTqisCvXdNeuQrhs/FK9WlICDJZjB+thaxA226aXsSHrqP8/drrU3BMOTLZ8iwK4bUY40DTZ
IArklULyh66NkLBmJYzP5Z2RfD8oEb1zxV9jrSrJ96EGIthMbWdZfES9LT7WNKx5yq03b3Gq23Od
z5zG6dfIZ36qchThORc47ztvzSb9vz9SEV70K5Lf536pcHiQbtjdHVUQygERfXa0HOWdpBGy/vf8
McP+TjoDXm8QSbEcXgICY7S4k2+ZICZe2wI6JYus891eWtKs5gClCNmtniQhZmeNPKouEUI4BeC8
yavTSCNlIzJwH4+sv0Xno4lE6+KQB+bm57tw6UPBjQLd3gVaYb9I78dnWIcwdXkCKe3gAL2mDdKv
1hBvrPnI7vPFwZYi2GLENQqJdtYIfhOWk0xc/FIaqZaKKbE/edChuSTkuUCt6KaijVbmgdNvZYXC
iTSu9yFCKdwOK/3i5xJRncOZ+O4iQLjxYFuQRbTS34JixIXEIuqqvhGAwEpRXBOOhSbUPqyMY1Oj
Yi0tuLrYzoboS6eRcfay6h994Su/Yog4Ae1aoQ4+A7qR4FnPa65G54VBgOXWQMgom2eWEDgyGbRc
AVkwxwD61Cw0+CNImw8dyTtd/TsNJDMfvDtF9yD2Gib6qK8JA1STay9ruCUe7CDRi8uYehv7lrXu
GZ9h6SZPgx9Rc4NRsW+lfp9TE5yRO63aV6yz1UjM+jQJaNUajz4r3TYym4TIIIn7ageVreIPTEd9
Dz55LlA6q0Q679+b4tKad8X4FEVF6+avIVMlFiUscbK6O0QGA39IXVJ9FSQbOk/MbSC5zL5dIeEe
xzgV2ULbOQekdu4elHHWQP4020T16PgbyIeY3gJUkmrx6Gjtyypb7fuRWJDE+SNG7lBwrVRM/3lK
TKP44MAKWLEDUqBH1prfoDkRoIYRCflpV4S9wJy9mMLIot2eOYxfz8hiR08HY3FaUOLCfla/hg0x
nMWBKiLuVf58BO+xSlup/u5AuaGEexRma1oEunarganQns61ww9JOEiomJVZcYQCXKiiXi+0+6Q6
1jsWUYgxo0Nxj4RtcIrzYDGzWqGd3KnhtlwneU2OtaKa+hxA+YEOvIls/rGMyONRFM2T3Luxk+Dh
w/JKWoqcsz2mazdyTKlTD5hDniVk1OSQDaCGWK0K6kR/0x6bkMVINSkeskNp893SSHy+A0E+/u51
qupQ/Gk78emqLGVT7NwtW1YeMRmbS4okFBzy+IF8L7PiRaW5kstqnP/EBGLJ1fpg4pv2yPCpJ2s3
/YSoYkCFPOwpz1Zc7ZxDsJmUUs2LqCtnQHIzRy5/jZaMXdMLZrLEOVgi6tJWheyDUDxR0F2DqBZt
3IGJPL44ac8Jr3zFY9p+p/eKUWlI403OfP739ytGawXoAbKrUiFzBNneQN9XRjLloyvqTjlLAf/n
0qkojeEjN35rYMew44eQ08xa9JGtNagzizgHZ0f9TPI3H7M3e5Wnq+CMd4LOeyJHHdbqtl2wQySv
KuBJ/iIAnP/n7EeWBPfVeYA0YVJ/dDXIOUbq7YoWHeKKr6zToCaE0SUwW1sDaAb1nOMTFPpOaEsA
PJ11+kARZjEj8uMqRoITtTWumTVkbeg+4e8KsYteQmOyvId+Y2aeL15CI15NN0h6UQ03LLrUKPzk
GzMzFEMQ5uSXrV+P78F5Z90RUd00amyKhzFQf5JRLa2kvG+h0/d3bSh/JGunJykpoaPTntkqi4yK
iJsLM1WaMm7TjkV8gqLdgS5BKrXzEFfLz1gjZwpbXIYl41qOVw3yMxLNupH44eNkvU5yWfjQ6nsT
5ZUQ3xDIYY0nec4qQ+FvToX9sOxIE4FeS/Zmxcw0npHOretVoHttN4yNPIK6+aU/vSYxihp6/6VX
E+5kVP7RprKKlNlVVZU5RYNVXgbdVxgtIbqkvjpfa+R74uXMVGLq3WXlrnqy+AIsXq8jkshld2d4
ghgZ8qIvn3nasWJrSTGvVuuUtKGzFfIe6LALfsWE/M/sQNIb8p5nVyuRpFhn8jFc7B3goV7TQfub
DC5doynoSAyYZe64yUuPkbIsekw3HtHO0EUPAG2eBNulcjNEv546DtmnZ+RBNKb2gKMfHoPDPAtY
evVdAMw15+0pbwRlA9xTi6x+N+DCXD4cXbyya7EpMy97xkPACcnnuOwscqfEMrpJiRJDlaF/cQyq
TS0Z8qe5ocGXDWLbN1qEnoWbvroxyI3hvJHVPs8HNDEmmlGSilF3XBA0hn21Ted2V5NsfMkzAcKr
84IzrqUxE0kssaz8mGk+y9WC/YzH5tkDRwWEIIonpT46q2rt7IbHPg+kppM4FIFAlz7RTe7+IQld
XKRAVkXs4Ysrapdgq2oxP48HVRHRJNRlkUJm4jy1hdk0tfaYro7M7HXPeicdSjbdnT/Y5zzG3+D1
1PNZE/TJyPMsorZC+wkcscxPLlu8TNRMPT6/d5OPJRd2YD/d2SHgAOmf3VCW7vhdiktboLVRsCmT
0mATk8oBvjgDe893v3QbpZQkCrMMfqOHm2MYTZFUMeMwN1C5eLmMJP/qIKQ8+NhdvBj06X2RCRDu
VT8PZCo1HnF3sP2VPtDdJW+UqOH4MCjLJgz3eJFSQukqmDWKt3inCcZTzq/GSmCWIHknD6ZAS4bi
pdmPEeDb1YO5oeXQLorxz/CKuEez4ld915S+SURjQIMTzlEihp+h4zb0YroEUJKqfW8dv6NEN5d/
ctZUIyAYhiYOb6KaAvLdSwjxbCypB4ejsxiKzVCJSfBjc4NYHJzYyxjqyWh8Om6eW9fKAYtA1RFA
IeE+AVf3kD7oKTHdSecUI0Zr0in3TTtn8BCRwfziqIev2cU9gyWJcn24zB93gRdeg6++8w0qlFTo
0LFzpqUUNMmjZqUUQfu3mJ0o/O7xUsXwJrSgeffxRT2XZCqDhzjUzpzEgaAJc4lETW1RAP3a1+Is
2tSsi/2607V0KpfDdMKlEK1OWznrk0GjFuZGnmdqF62m9KD5r5xED2wL1ZBPynWZ2yinmBlROHBx
R9py+uQk7EDueNl+SjjxD+KHvZarbS15182K60FwZ7vUwPmIjQdQe7fOtuSDCaX88t1Mdy+3PdrA
15BXlLI2lhllOhNhE2pn/+iWk6QsL9o2/+2hZt35pLwSdeI1wlZNWnZr41eGChtrUUZUUTLMliOC
6C0x6Cc1sxWOFc7v+NFCe/6NG9nLtLfWD3gw0zpPB3T77AqzZKXhL9wImdErcAQ1k2n2cMBDSEYI
YYf7i3ICIA2SdznDHkFd9dH6yKCS79VNxjocXCy8x9WR1AnOs4QkCB79/bq/dHm/OO6Dxhy25l4X
OViPK29ml2vYj7ywSCja/qPnrGf1xno6tmazTR2gv4ZyV9LmTLcfzy1+/iC7hIw54+T4vAymrVio
u4lVLmZnWBuBC5WvpNdZJMOOvD2x3qaQbhagxONPDExaZBhPcL2NNcN1hCBYSex0AbWqY5gtVTqA
z0jLRD6fzc50OyeBOylpag/V6Mb3UshRji+g/F4HGbxfaqKHD1HWqLWdb1JqFP7ceTAxTHHRpD/E
GTnyKMMH78rWtuwpotSFDcRmDDcP9CLVs9oBukW9nN/g1/ZvICGx/KNT2Pc0g1JxRp+FSq3SIb1U
wkJZqq4DiLEfXKuhvkhgoD4+AXuYS9dIgIFgfQbjpY+i+GyVz4A3BilFes+64tZZtAo54266RW7z
DjVTFmfJKHku9VFDWD1xCQBH8Jw475gavDa/ZJvleq/0MdWhXISoIpv0EtHEjThiZRnyXBZ4aVvW
sqkhymQQJoHafspiRp+IlW/21UEegAEIkrTbj5SKrwTYNBqN2DkGv5E1BDDv0sv4IzfjBFIH2t8F
TtZFEztEY7Ni402ZxDPj3nlgf1XrXHETucjRmisnLw5K8/gDyFBntsRQr5NZ4uDZfnmDtg9lIJC+
t0D9tW2r1gFXKXV7p67AZHPnWVnvbzcERvKd+oju0QU/O7O73tpqaORu+zQs3GcEmY1gNxvTOpfX
/iNcOTdypJx0Lqdjv6ohkABDeqjYFx5XCW4Ca8W5N9LRdeHOXmewitH8Eu5sE5jQKauGxhTAIS4Y
MN7EyfiJDjbTZ2QdxCjSU8uV9KaFlm44U90gSUaw1prMJIf8kQpNaKPiORC/Pc7ZXt3GgwR+6G6f
Y+DbndpLVyndt4MWSy1e/O+MLWEsIMkfOm5r5yKA8J8IGgbJKq4k5zqiCE4bgbp2HEsH0SewXYwL
tgPzkXQy6cJ2N51OZrKXPPwQXKCCsVfOEYne5flQsUQ8c0kO11aCJFxhDlmEIc0LkqY7zEEmlf6N
72FoIiBncNIoyMX5AZ92HOzq0wV5qKHl9BMNp1WnXPVet1tdtxiNdcz5vwVBsvD4PlkTeud0W2uh
oyXfx3obHNRvFvI6wcNCQBpn87rnRe/d34q4dpUtN3qZm1ba5DQoVlLaPNn6awpkC2FDF/AWfKhl
A6UFC9pok6sc/yCyYlQhYlhkWH6XmqHlv7jJsZ3gINA51PRRV8pOummJsa1HMwd1wXEjBBvyWQd7
mT1ym1vQBzXanXm3ND4WvP16vg7ucV5TZRGi7mZUh4vKiJV7bi6RUkG5BjhDjWp5r4XK/NjAxoER
jpHIWvx65WumlygMUo7TLjsEfm/wSKhFCKOAzkTcQiG9JNG49ZZKLRbKYO+6SdWmYgltR6gO/cD8
EF8bnnGgpQc34dYsFLqVlj7WNiGumAw530JT7hP2WxaF+8QrSKFw9JFXPjHDAwc+YNST/IANeNP+
qrLxoClhuPD0SNHPJDpuFpxFUxgw74oyuU+GCUFKAWszktk/OB7M+Mkz1NAF0LxnBFGugq0b5XZx
AMWhDrPmmv7W0RWMPooy9zE6nzddSMN865oF1y5BsEqWDo3dKJD7pGzdWee0WJopNGBmBc+eAZNl
rum9W2yDft0UsO9QQQKpFMMN7ohHhYqZOEUTVnmipWY7jtp8Y7f6eUktwBzMbRdDlRzVok2xBOU0
ghQyPy873NM73XednBNsnYHnbqVYb/HQQ8/efAYsKy+A9fjfUEXH2DcXh4degCjtYNupJwJkXI7Q
n3dUJ1FT0ul7QcsSYoDQxA/NPul75ViXcw69zLzk53rVC7qYEbvnoyZ2yUiG8bII5OSan5zp+uKg
HaLAv6dULFDGOWEmQi4bw/OAfY9kLp9C+09yXZYX2ynhumxvWFhwVbzHFWhOGMfXF2P9nsbqa+As
64VUIa/VcjGfIzVXdpbu79evS03SCO4cpQ8CAxASkfHE78orZBGaK4cy/YCOOyIxFislGo5lNRUw
NtVhXM0CrxdooU7u9kVORLWDFUAYJKTuj2+RXT6eh011klzlEs/B7+3tonDjVQOMUBjgQmzx1d/2
5PS9QunrzMU9GKWum9TbMaSNnd2P+fpoJMlsmL+FPDdoicfklXufrKzEfh+Qxsu68jsHM2KdISmj
9KJAGua7HfGHWpcgLxBDeP0v5uRoIS44j2vOAO5utHap2sHX5QHksI9aWzR8/CPjgDOFb12ikx2F
/aTvEiUqVbMZKDJBWeZmAPuf6roW+rPXiyIIjGhmx3jEWhmcLWGWfdrlxVpwgtH+UP9oyU9jHLBT
5MPKkcH88BbFaZTymeiLHDt31Uywp56D0XvfqearQh5mfglLYUD06h7rYwzxRZhuJzDH8gPJFHyg
OMkI00YFcxISKT2ZRyw7N85jsCMKBbsrT1UttoXfGuBq9uVftbL4T5jjdHX1zKmB2TIn/lQPYeid
JDUCdHLdyINTcFDtweorgxy4PmZw5co4wR5TZEeDtLqscTc4VRzz2DAaBQw2iS6LgBW7NzuUSytV
3qUOX3Gsfwkkl02TmopvH6i+BZp6ejdSUDQEBPC0PenLBukso/XdRoE59mFBDx/IpXsrk0zHgosR
WXxNfJxb3NrwaE6qAIojgjvtycbF2gF9QBmKwxayorcuML3OXliLv9WC3e32xz1BasB1lbJaLRPy
xVSlVBkqbSZbDP4qprexN12IqXFpBllEr4A6TaXZNxQgXSMm++XsxD7ohKtmC2eoEqgOi0fqyL0I
v9+luQqGSIkFMGg+5zA4dO5i+OEVabieHEEyb/WRWg9EhjFynHHOuXeEyzWZAIc6zv0g6RD/Ug4u
Qen9OKHqIjbh1Uwos7NYArV9JM025jIig8gtAX0o/ecMWqZU66S0sjpGkYUbTjeWvqTSwsOXCWgW
y6HJt0Hs8Kea1DGy9oEuOSYO9nRaECkBuhH33PzrkE3BHvzEZaF6E89pO5WCd4YghWYOL+NfE0vg
XLw9UVMK3HNiLMh0DYOaAxiGRGnRPt6luFLXHworQt/HDUyC6IhhJJr14/TNphkvGP15cxX4IHgg
2xqx498SPPL8u9u7R7XdHp3b2ggTMMKisQLcAtYgYMbRgbPe95W5G4JVXbQjbjhvPWKmezr800Ps
bLZ0ncX7rCtLslg9zuuCzm5EPLfvxmtYn5zSmlAMi3wWpZp6oKxPQuQ+5PBzrdBJ7G2iLAtdVFmL
3XIaE7Xya+yNBjFpNGfm7YVDNSfoUd6T32qXaioyNcx8USNikbCU/RobrvOJX0ALEV0wwDZqKn88
/Ply37PufY+Elqfa+T65b6V+9g91unZtZ2DIP+MDi91fN1qzWERaLHCUIT8jOo6usTj+tX3Y0a/6
u3NkOEC1hWEadoTnx92m4LoguRMauzlVpfKSJ8r4fQWycoqwQVx4bl28gqDgJ7fNW4614vPwpGkN
eQ2O8Cn0iCEQlmRjPxp6aXIMar4cgRNK8xNge8LbDitEjjXvaBz6EzFNeyGK/uIjf3Ht9ZQryhaw
lInzSgunheky3o+rmMWr07Dd+1xIUZLeqMhdJb54bMfqm87YYb9eYZm8jr6118UHiEYA43GgKOwR
FbXx/e9OTuxtXt7Kj8RqOTPNBLQ4wjP0QIYW6bC8acUX65iKHhN5hOH3M92l1Ph38ssbljl1sH4J
5fl8k+y0sxQ9vNoHj3/gu5So/P4DFZsXlFbnSfeRsUvNTfkGKA1IBFp5VMsQJO2Q9ZgKQsRQq9LI
cdluH2Ntl5Wu+usDObEQz031nUllIKpWz2dDBxgDokuk5BQS9uoAA0C2LeS3WAxNuuD2eSpnWiR/
kzdsF53VHq5LYT+rlynUaZD7QHB+mW6GetUXNV5MaDXkx4irRCK/gIV+dUItP5rl1ZXfkZ/+bGNC
3csOYwC99oVRDV5Ua4NHc3uBw+zJc49nysiDS2GUqgC7Z7a2rA67Zn0IbBGtyBSLVe76JBRUzMPH
6REleyNFfl+oICfP1dK9iFdFuWMC75HuBLMaQe5MQSzj5AhUCstav/OGm77Z0/NfVX5MB+kX1mmk
dqNpNVwlMGS7bA2PRWsdbBQ3VpBjzoc1vs3H+3+XrFlkmEiIq1gGbkSOivfHreczeIUIbgjYxVNi
7CyqGWQ6YpOF6N9UgJHzJC8wlfSf5WKFDUrcQ2ZYRqs9VlPvPoqr7sHUTEe5y5+CHxlKIFh/gZ8U
gRIwYbtMMfN6XFAZeAv/Ypo5RKckbiTzHakWURU2wfOqD4ZxoMLsfQP39ug3gVYlpK0IB234Q7NX
0luX3RxV0l0QwVweQ92tZFOSCHrO5Ox+y8DMtO0ktsFu3Ukhx5pkWGHwLKddL87cG7h5GXxkIep5
X5UckuCUaGThJ+SofAqRjLeLKlcjoWFzAgrRLrqz09kKHQW1Zi4Arfk8WtKblLPHrXDzj41ETp0I
Sn4mBd6btWy2ImxcieikRBtq4ld+CwskdHctCeAl4BXD4UMAmF8d/iCaXqDOv/4mG59erpsGDp/a
vm9Efyr4cBdqeoTLMfFTDDZA6E2cZOsUZGGMjT4d0Ro4X449dI3wYAZkt0k860DFigfgebrX+d2F
ojv9yN8fGvR0kUJYqQ/9UVPAMsSTGEg9o8aH3GZSI9k34s1VDF4xlQzLvDqHNrHU6Z4wDNzTwGUb
oUIqqovXObroij2fBAQVyJICsuMaS3AZdy5zAGs6Jes89F/hDysScb6f8aVfRBIZfyiN+hrYg6Bu
jHm6g1oWQygYTDxxQYc2dfd+I7kd8S7F8C6Tac1E5BW5DidSa2vqcucjDT9QOCBclbcqsvBou77P
pMTb/KefOpU0sdKkVUBp1pNPjQzFAWxU6IeHsEOdyrL6+LYQCi/Lwg3jrzKQhKHEjW4X4afe4bsy
R8GLhTR311uihQN38kB3cJHUeZrfHP64Omgbk6KzLCnHG4+Sm5jOHFmkAQG35lqWHYZk0eLX4hyF
fDQ4WD6NvD6KcrwzAkZruqqNKsvPET8zAnFEG5eWE+B84/2YXNcWVRJhcY/h9SAvbQQHuCmRzlJY
tZnqUktEbrdWCcomlxHiekCtSV+geV1sPm8W30pOch40l7HjsHgkyOBskWFYxpYfBiT0FYs9QpEf
yjXCgarBDvKE6LSxXav6zKSJc5ajzO7YsSVt0FrbPSy93BdqxZVGzWIZzonlDzqPQ9dD7bQNFwpK
YZ779X2BUInZfkngeR+8x1WcmqyPWre4G4NhvcDuTaYY2+WBej3sBJ+YuXtLYUAIFSlvJlizLXsV
gEUqdIc57PNKfvoe5J/4ptQS2Bg/LgWZ94oaLJwyqz5kh/K4Al0/ZYGozlT4t1g/jfdbCHAMQHoY
p2L/S/aDV0Gcb5vG0fu1RNeWO3wpA0gGvx/7HNw+XTHOlkgjL9/BSGYFZJhkmw6FCNx/CTspnnp6
yvZfvCQ4GjgvNJux4GwfVLfiV3mFVnH1pzV0lycIslHb0RXS4QEevdFdUgUzMqFOHpo4D32k/xSd
90dZ8/aluyzQtyB8gMdCHxybcnc6wY4bLz7FS1B4AhYCLDL38rW+nopOynA5PvXALLQxaJCx6Uwe
hUbwMZhmMwjUGYU9drgGHN8LildH7mtM6SXTHJ4WPX+KaYyPWsrMshooQPQNZDOVezuiS1y9rHlm
QT2EgkSQzCnmchPzQ6h1R4IdlaHf2ypDTRrYKFHQlZpbKmLdck8DkwobHWrpXHt4EGrrx/HJdqF4
f/gFgd3SuHO2MM3PzM1uiCBcz9CVkkD5l+0lnPJfyY++dnDNFN8d5cioYK4AF/pdZAeaG1EEc8fs
iyP9N3xiLNJT1ecuGtLGfUlQxbeRHZziKGJQq5wWDVmA50unDuU2XLlDrymJMv4sepJEeDYq8QwT
/QaBYFGdiy1rlDrb+l88n9kUdtrv1sdHZuof8+fpdXocxxKCNO0ag2O0OsGkSzn147LAi3pPTr8F
EwGaskA5E6rF1Oc464KY+CY0gMPFxY5fns2fw4FzZdxRM+vJgpK5gmJOHDtD2rPhhgEjq/Ycp4bX
QbacTgmRrF6GTIY5DWplA6oyLILdr6TvH3KJQqs2O7Joa0pfr61HAdc3tHu5o0fQmaiPAn1Z0fxI
/C6DOZi2EXFstqcIKMb+E4T8bgahacjgMz2VE39kyfNcy5AKOfKloNqKzcP3VUJ5PxVSEBmDalY3
GnpvofhoPI30QTaDFhlX4ILmjtUGMO8HujOqvbbZvOXXeoyYY/ZwsIi9ngQYd00ia9jB0zPY0Lho
g47ce92qauOJkJ/3yisC17yqupm7MEBheG6BgLYcblO4Rdxkyb18nbU/DRjXNZy+KK08N7nv7M7X
/PYujzyFSuwOY7s/eEnIuBQkha4EF8+djnF6r/zolUeyqaRYi+1xh6T31o+Y3wqQgpnUyJWP4sKZ
rJDH1MGEPdvjk6vBLzup7z6oLH3vO5rc3cV1SAbwDqt3bS+vXeak3ERydXb+2bJPEdX6FmLnA7i4
XbBqzo2tRLTYDTHYAXvoG23z0EteE5AQktG6kNMPsq/GkIO6MBkjiPnvmbEzMDWw9zcyUbhhH2Dx
FhbrAvKldDJApI/67MQoKoCBgaWeN3gslLcBzdU1fX0StsoTQc0zFKiJmHRttTObShJ/H6p3lDYF
48UYKE9N0QdYjKlfbvJ9y/QRlkmV844MvWt7Oso4kWbuIjEuaU8PqzfEU5U5iND50aRBQya3XNwd
RwqB9qOlojXJ9GB/NrzrBTnqMQTMHqHYOvCGhjHJ5EvmAkJIl9KYqSVgoRF2E4FuLGWPqlgdU4QK
Cx6ovYJx6flFIXsLSZdRnK6zpoHciUx1397m6NdLzc2H0ye3bQo0ODR1Kl9d3hTbTqKJgrqiVkyb
EVvKxf0+4fw2IFxFrYgUuvslHfnentEeA3nEzwdXI4V/78OFiM107MLDzMIn91agXuAbsaXo9+BE
+gqiMTHoHEPI58AYL7Y/GXftnGXjnnA3/f0/caHufjibar6TDaDm33UUn1EsGazkrHaTexanoKYC
FL4IPJ6NoLiueb0nTQ7pdnJH8v3MT4BQYlHJyIL9GZWkA9v9U2mdLkAaXc8bLIT6GtFlHHldd0x7
fNGza4oNmaHqeqeB33LO1V8UFJS4/ePDbuoQc+nnT2k2QJwAMhTxafDiwgVipmX81hoXLS/tMyQX
DWYrIHH2VEPcTX+gQTBCJ5OHKJlTz3uOruhbn7pTKukPwAL/n5GKGqlLiFmXXvmwSXlPZ3QmXzHW
zP8ujQ3yJzSbKTIWvxcn21GBX2TNMlDxGP7PYRGSuPMV8Kp6WTTVziR4t3z2HYGbfqqnUfNDzhj+
URHaWdamEUDYq3R9E1//s+Sb2QYuwSNo7HJyxDIDvk9kq8fY07YEvI2VWlP9DfES3S6P0ZlJGnPr
vnIFycHzeQ18Y4cgWn9ArI5TbIac1ssCdAJp1/VR7r4aUJpNYZhlaDGdKlGGFfBjdfAftTMayArQ
Aceh/7iZlbHVM+SN+eZY+TWd0OzF77gm6N9OXfz4aUUOFWW5Nb+LU8SdjV/Do2womn89h7/3vAIh
J5al15oLk6sAmCSTjHGRJpiazyPCUbL3ElBIhM1SxVGizwFrkPOnKWLvxCBOIllI+8FV3bdmTFf5
v/ouviCUt+6k9SQWaBi/02tEi9inxbWxD9ithjIWuluUh2QD3L8HBhTxEJX8ivPn8DAr6Nrx7NEK
UPbyUVU6Gm1e07xpp1oyYWFvrpJHJj9GGpVI/l4ntQ3Y16fslDhyKgEJrQsCGXaY1NJQc3QzUiNj
LjCx7EQ+scX2xweYjbUqfO+DAd4Nc/fqH9p2qOA5COfW5zni2FpMA/gxoPz4ngkwr5fywm1JdH30
994fi0vazbO6qXUwZmCvwDvyUb4ogX9dUmjCdiSfgTa2B8fgGq+7LV1x4XCw/kzR4DjIvrY2SdIA
yhkUNdkgghd1iV9uWSmGmwjUwSridqfofcA/VUeZ/XZ3oJmAKVBOQIcVQxwnAqSwNpZJeKOV2im3
2/gWeuYVFawcSzJs6gHpohKAfdRC/pteW0pXHiJ1zzSvv+OJzHpqzLNxY+2d8DpNg1Rwpotoc3Z9
xscNMKVfQzB5p/BhM9GjYSxIeBWQug+vCRpgWhUsjLyo47S3uVxn/tuF1cG9RbgTOTd8OFaTn3Kn
g+yqjiZmMJGKmcEiEek2AITFn9RTx3jdozP/Z6GCQW9SlinkyYM18Dxobv2VxaHsVAPzMKzzUL4M
ZA7uCGDWpOqj03hewXHtNxKMcrfdWM+mc7rvdLeQMTA0MwmC/02JWvvGahUA9gi1N8b+tGC+Prrl
42/bfCODRbDBzMMf2Z0syFXoTWI7r0Bg/hA9CYhb14k2OLU8BPDxnDELgJdTqVf4zM9uGcFzWnjl
1M7Sq0NoOorP2+QmmumThvpEqbtQAK+ZhWIHSUYVeE4qvGS5Irf785RIr8NhyfVTS1elbLzwJZ0N
0IR2zaG2AOGq5cxQyZKBIKH0irDGa8iTP+qg5uL+gdWVfPpLaE9R4rIKaNVWNkDGaDNxtAImHPKL
b9+HBV7N96A9IwLYkVkpD5hT8ibmWO8qHJZmlje1HPYR35yMeJTOgy3gmeCh5MMjT76NFOrM5SY2
qB55XC0NCYqLdSeX6HiLcvWYho8ior7trT8N1M9fdzbdXUH8pO1wwL0DNW2Itmq6dpQ2tLsIZz7J
BcvKyuyAhfyghfPUNu1VwzPlFEn4MpfYbwbsSEiDuM/wazW213S1SONDJ7P0GxAgOt6Dxn1+RQMR
zS2bpj2B9wePr6Ymcx0OiWH9gaCTCmN2/P9hLwNT5E+vlGUhHJSdZt8PocxqX945KN36fu/S+eFs
/Nt+S/YoBKSTs6/fbEmA4ewQ1TsKvpFQ3y6w3OmdibynDfmuKyGFm4UrKARbWmzN/Ccw1ZfgZUVH
X6O5inc0AKdUTUo3NC17jS6zkYaqksVsdERBBhx8v6IOjBSEPnEmYyOaAs4E4zt2/mpmIBHWk2uz
D35V5J4OGF091m/qlVCn7QNjtQdg6k+8HGBWcPRaIl9WGFiMoiFPgH/q2KK028st0G5HQakzznlI
TE3EfOQE6dqc1TwiPTP5e7ycCJtHUkbLs28d9MTT4ulxcZjNVS3lSEpcET3POAyWrtu3TEyQ2paE
6zxOuiqMT1wopLIJn/b6lfZRtrriHWtfQ9mtir5Zo93KEIimfCfhfc3XItKRuQS9YfNKKUeJHDcD
Fj8a/IZCAgja1WMyhjc1HYlku99W3oH0MGT4OqDHmfdaTvxRTxWRszQZyFCXYJqg+vmPoVij+l2o
vSuZHBhzh6e+lkrlqadWtnhrsm6pI7eKU1UUUlBuTCASHUCUY8BL/HF8vv6APbVDxjJ3WHbHrVDx
BXAw36qHNQiD5r+CQjUX6YDujdHcSe4Cvg2N0M/rZeSTLAxd7EdKM1FsjLFYajnja5Qc0MBjZ7x2
PFlN7+twx608LlIwj6cpEnrQADUL5Mo6SunYGQ5bhfAf8C0dM6wbhAty8+1sA+GvyiLe7LIiiE9W
E5Nj5UXLhCylxVobixmFfG2idwXo3SqBwJyQJ6Ca4F6+XBpF9FN9Nv8HMhRe07tDpXWL/1OrAJ7a
k67eDA75tPrBb6mQoSrZWrLpnXbCNh2mQCuPd1umk1lSrePvOkpk4gg3rXwduSh3vtKUjPOvvQ2c
V9NOsFIXB2ZdEkpgbxqWEa8cgU4lRH8xAgTj2VTwATdLxpdJUHXUKlBBAQcQFS+X674IuZUkyzhQ
RWIgqBobOLzATzyGsbkZj+jT99s3Nv3Y1RrXEJckM1f10+uit14o9b6GHTF8m1zDw7vsrXwJH4eT
/kjB8SE1dCR+ZZzREPa6l/nO6BeXNkE17nHhe3SjOX6cx4dXCxIdux4X+jk/nhekeeR4nNe8dJeO
yYY5XeZpivCpkU+/KPUDZjZwfQuG0fTLFWxmSeqMfPrV+db6qDYHxLIpjCGT8FdgtwYxgNQi+V1q
e+PWE9AjEMLw9Pr1N7w1uWENTUE9y1LY+LIM47wFDV8ohdr4vmFdGOG5tKvmKbpEeFT0kt1jH/5m
kEG/JkUG3MbLs2jkYeLzOpZ4ocygnKHftPoGXbwS3PbeqJCdyRz0Lteie3M0Zk65LT8IdhpUfPU2
kRo6qKhUk2qa2rR0EeydnzyPwflmJVljDIfEAtgaJr3EGiYdK5j2eBEio0Fe6fZVKum1rQcfidHi
xYZ3dcvtM9It3JPUisWJZPcvHJkGB8viYpDme5uzp75zDWPBOGzcA74p9BePJunOkdVF2Rud+Grn
zcnQzElWQ8lcQRGDAbKZkUCoPH8Rsz5s6hxCemBX+VV9O6lu50Y/EPX5EO9V+qMSu7/5M9eRBk5S
QAjPJCUswQ11uW0JWEHwEv4dF3vjRxdzMXqtRqeQ2GK1IZZ5+dw1r2k/0NzxR8/E9UMplM0RA1wJ
d5yLYJ4qq0LTS/rmNRiAfQqF9Zr4nDTNawJ2bOxUy6G4tfmox3gIEKfDBx4exJMp8gGuXcZs1/Fd
i2n5BzQuE0GbF61p7RqHkUA+3n2J3fQ0g8+3BhKMUjRNnmemtO10tQqO8HN/Qrzfhu1H0qeINp6O
0kI8HQhQCDUTdN+PFdfdo4m+9Zg7BLVX9MpYRADAOfl74svNrGklpWt+VN/2XCuUuOq82EgHVkvv
S2DaaovIEw4Lx+tJJ2qLTijZnVznxanUI1wRK8jkfzSYJJMw2Y3CwemRMM5SGXzCsUA1+RNTEFFc
fHDHJIhslWzIvSgFQ2WuMHyZvRN6G078NOV0cPO0HHXeh1oyzaw4JxarJZJ8cT0wpgpxzZao19ii
0mlYNHi5TS5G4a39SbvVBConeDzrwUwjMUnx93dNFG+YfAsqsn99tmkL4z+fqOJAvMzXAq+1+0Ou
8N8U7uaaQ939HQu7cnp3N6Nt8i5lUsnK/3qUor5S814sssHlbD7IPl2UPkPfUoWqtyKfath92Y1+
8Vr4zR+yScOfnCvL6ITAQvM+0g1FdMxn8AJB7HIOZScjy1CS+z0oc1jNFrV3o3PqoQOjjrbsn7M9
pICT0ErtlbYrdghYk+i/ObvlpqO7MaZutFQ+MQw8L8AgYNyfBgqkpyzwnMwd6JeoVSz/w4pHdol9
mxuLHAnvcOQjsLihbgFNoUxbEKII7js1KmOJ8BDsh+WbELxiA0JjiaYRmDUaM0IXTwOJTEjxjkWP
GE4cuy2LKRQCWSTzlz8qEdaZVQBSZU5/4HBPBtcHy6TJyZYk3+sMjDaJhO7ObvsYKV5PaUzYBnVk
lUO/pLN5Pxn0M8WRBc1sB/NqVx0ymNPKsYEXX0qBXWutNEHWgj1Ifz1ibeu0gHdERveUzDL0OVbm
7HpspGhV4CR/3R2UHr7/cJLbtTq8wKyUhT0d/+7/KQDfA3PO4iZ5Kk7OxymEHsvkmikq6BP8uMcx
WrwFXXeBpN93cAviep2XH58XF4Eghbhf6blPcwO8EUERJJ6c9ZxS/MbqOhOfFBwIeiZaq7Hp7czT
ZGuTSBkoSRrt3a7btBbV7yxp34PftLxd8UnorVu43tR4vLIb0ia3K4BIIxN+9JNZD+lfTr973mxM
ay0Y8fIwhMvy3hD2O2duPghzFxFYf8yPapmJlqjeREePrH0djDo1BfDiktJRPebsmlaWo8zirra3
XalNDnXRCxi/KmVqUv+zN3/WjeK0sKqoAeJ17iS5TV9SfkyMuwvMv10tiqSvIRcolxVzf6w9imA3
Abjzr+OqJpxdl/vhHYiaDkx0m9ijaPWlv3J7Q9WQcmH8iio9QNwUhdZL117fXs1sTfjKCZQ9EiW9
ti0N7LrEz36DdPzeW1ul28tAR64sq+wmDBOluI3jzGAceNYaLY6hTI2WJ+OqFUSg2YFt7a8Ez1ja
/zVFmfaz7ItuKRH5sf9jt/PD+oh1l1QCO/32CzI9TKDpLxlgQyjPRolpt/iWl0Oll4QvMgC7SKjk
WDwCeljeEqfygIx3+Vuqw3r9Taun5VDp12rX5OPnq8vS/qM84EkMmp/iWTKPcgfILMyejx4GcaA7
x7/nTX/KmvygAN9wC9xjaUDxe6OGbWQjjpmcL9epBHZBLfFED0kSZoCi1EhskgjssXOHxKoaZ/Wn
Ev4Mt2Blj+7dlqbY//g/c4NHx3MCzVEjG/emh+n5wYmM82+gVEGQmGVq1Aj9Q7fmW4SZ984NVr/2
92i27J92go7iHUuAQwFJ6qbSrfOoSO3an5/H0cVxv5dAQD4eDJ7C4tSAetox3+OPGiH5qsq0ppU0
AdasSg9ENs5LQP0msCSXRPsTbUg9rCPKOu7Is0rnqMQspWS5h/tOLSVGYALKd1Rs8KPt8S3rBzMy
mhgPh/q2r3l465xLpf0f6h9tY9Uap/0a+UBWUmiKxq50Dty+vp8ayWTr8YJ716QxDftFSqxfomdR
/Yw2YWsylsFiOAqIrsAbWJgO8LR8QhIYtALhezgRio+GV/+Gh7CANRfQuRhRXn3kH3LIx9+h8JLb
JsBIrGL7vt6sbnTZQXr5UsZ7UxN83hvLtY+7xwscVSg4PwrfmAJ3zkBoVAlVLXNbltTlmGqF0amu
JDs4HTDVUf1ygqTCCzAy15UlHTgjUjjZdtQNTmmU63HdU7XD31dNtzi2IQZsseLG8W9cUEsDJL4g
xEFdTRLCNM1hc4jaUacRUuFVllIZ1c2jLieiUSdCz92DwiPjssQBCryyAqocv1gL0Dw2eiOYbfnq
0O/qzlOcsPT7Wg0be4+IUahYIkWaPAVzm5/W2knc1qfC8nPfV19emmIaPP6fOorWTrAYXxDBIuL/
SiXX1/d6Ht5Ie8Ji4xWtBLG4oVQogrdurcDgn95J1StzcqB/KmVPxTDGZzfLwrlRLZNlpZWOhqXj
X6DjJwAYEJCf5NbHJS/sT6/WbrKSd8kHJ64XE1m37cd7mAWJBXNNMdjYDyseXQwK7Lw+1T2GAmoY
xP9g9StCeN8zUupDvzVGQdIdj6cEAzxt+derJ5YB3a/2dg3aZ0PemKB3dQPUbQVgeERhHCb4+dVc
lysIXXR/gbZIf2faHH4t7dyvPIQol0qQEsFraZs8CEpNNvNtL3c0RCfl+svICucU14ZdesxUB/yh
jrUEykwXZvi/QwYYclugqq4GwJkbrTQxRQ8EUh3GHs7l6zkYnqqpR9wOolUBPLD6KN396qYuE5z9
5ocScIGkieZhyDZ4wNlRWFO0dhBlvIsoeqiBVAA/1f7KkmcRvuxDVZKTpybJBdeKDJwXFsiYbBcZ
FX7LHUbegvAIG4df4NV4N177DNJbKnakKk/WpNt2gGnzBa/UVUms5eP9xeFe9IBhMZMuS8kFE8/Q
6f9tizzKlm6OvRYWZmqzGb+okOPIEHIyB5lQ/m9mRADEKjmj6yhOV7QJ69Cbi116NsdVt0qgnPHT
ThHEJYo0sF3yay5UZqT6TgidzhYgQwvUc7d0Ea+FzbWq9fM0yVYGqZo5oYpk4uxSbYZCK5Z0Knmj
Yj6iaCxMHbk1Kzk74gKCTsWBxSCO9ms/SbhhhfASXdOydPXaJC6w8fSx5d25nVa2blxFF+7ezELa
ZoaQo6gcYQEO9R2ILOGKL9xoTI6oR/f10JOXL8IYRp68iLtLtx7qMLi5VFkz6WsfOG6vkfqb3l9N
m3IqaLuHB00UCjAByoNP+JOFUAqa/x7wfPc1LT6pmexiNSwv+aySrPDnhjZ67sMhrL48UqBMRKie
T7shMc3pN+eRK/p65EWC9Sbi1abbt/NOcPVX+bhzKnikrpwBzuhiPgtE5jmiXcwJSa8qPVg+YutH
ySvEM0iwvi6uI0055+UqBNTmg8RqnIemMFfB4En9qzoQ7pNYDKBS6v9yWbNed7IwM+WslgXMD7ap
LRmMuAiP4b3IqkNgpZocxArQarySvb2DrbSM6imwWPFDBXc8P8fklcvT4Lb0jkuMK6y4JNu9MiPT
gYak+Ne1eh01RUDm2SEW9UjKSJCbfLpkicDMwKBWDiPKAEGy6tb9vPVppQpA1S5+rHNu8K60Gf+7
SZawIIpIGnRyKxf14K5JDkurAkfT8s2TDYq2WSajX1HDPNXyNMwwzB2PI99cxKmRVDfmqU3pbqO2
HjvZ26u9JrAyU3lzxd6sSemPBS8sOK55W375r2bpXMhIWIITQabc7mIKLaVAauiSitTPcaNRi4Uz
QxsnZRIyf8isXr9urPT7bXxeY43DKLqdNMkwQ8RvbtQJpAM0iwh27oC7mB7/nA5EKlV8VOc6d3G6
Wgo/cU2DdaZShgMpmPmxpheCV416EbfhWTECCZfhznErRyQb9j8Uh6x6KobqYz8LiAqETeX3iVNe
fR7IE9We5XLt3n2z2i+FXMXF2vdp8w/sNB68BRCRiMOHtJBLJqO62Bkwsr055lm7j5bfE4esthhk
fCF2h662wa9RsbCoa9OkwJmnN0P/6EYdg5SWBfewcUmKysCeLouz6MILn1FvZtpyHkH2S/dggv5d
A+zDRkxdXScu87YhCypQOfQ32n/tMEzrEHmvK9zRBUAtoYk69fwgpaf53qoJaxq5ORKM/2KxWMKM
dRahThfYqveLWSIfg/8unqSiwUY02ZCUvjjYdDNaQi5AXDz7uqs/2Us+nwlM9w/lh+YqJcbrqMSv
5S3pe2/NPK4cHHFamrH/r+Ucse5KtFhgiFBov4vnf7txwCK/8KCPkqmCfC8i0uCFkhlS2+KAn0dk
OWm6GfGM0jMbHfYvHPdVFoTqvRng0t3jzqXwnGY08ENAo15dg05Tq0ZnY6ifP/1rhuFa54IaKit8
osc2ValZQ99X0oBRAgg8gzIdC0RzanRQKsu/Xrs7QyrTbordaCahsG3r5WRwruvhXettv/6cpfXV
eH+QukBTCpcnLb8qZOc12trHiVrryAnusDQFD40ZuQBUcs2ejbUTIp6JcENJyShWIGMvAlt5xEcf
6kHa1e48vaNHha3+Au7BK2FwDMFusMWrJjP2AgKHnDSLNBjAOlxBHw79Tvgh+P+DMdFEgyghgigW
vKF6TksGlJxStzFvkWZWJrcNQ9AvkU8j1v5wad7L04t3oTA9HF5fWknA7aGhSE1Z0ouCgVMugUZU
715v0t+YbpNrnHjElhA72+8k+8FZMTFlkEx38849VhJ2zVzbK51QAfv45GowWGALs2zi8zlE+XT1
6rTAtptQOPCWy9PzJaTr0nYmt6Dor/fsr+iUZnxHUxV0KHx/roOdu21QtTSO+LZUNypwKc9glg3q
4UZx+twixkPCoku4wRCDTHXEPuEJ1ILEEn7vIxyPSloMzng01LX8rhFpDdvX+mMPiErxyzRgGidQ
u9mtebeGxYWDtZrFViUdOftUwXxfrpv5y4pbzfx5z3BoPXeGfJRZSigmLp6+I8mlzgqQKw5G7P6X
PwYYwrsKKXomv7VZ/UzesylyH1+74Xl3wd/K/7hEubATRA/ntoYj4pmoFXJQ9V5G1velnNOma0uB
yFNC4UovhsaaOjWvIZ1YhGJ8yKqgyvZLqKuwH8w/4rWNmhklNboJUmWSzkMUy/Rs5aK79N87RsBr
cV+bcLxRp6aIaEhU4WI5mJL+MYRwsvqM+7dSYN787zDL4R6OEIHq5Id+AETJ0F8CHk2VXhPuST+w
qEJp4qi9DG/qlbNnHtHqURRctXnRu/YJWw4fAPUsI0D0UH2CUTmB5StfEfU7C45wub0GxF6i5YvB
3a2wniC8zx8yfGax/fU7A9LrKCbzkNWvDH4eizf50X2tUkQr7FJLwQUBoI9CB9kGMAVRr8BgvSxB
rtZBpfkPIR3Tz13DxF2++D/rtlRCpG8e1FVuuh708fhSMYZIhnioLjiOFBt+jRf8mM5tkBQJ+MMQ
A2gRgkgGOGPWE9hdsxhe4pZ8P9qz/MYrtuAQdDQmpqVaLXWSvraxZhduLEQDP2I6TD28zYfFnhzJ
7jFIUmvoXbpKJdJeGkJPVJRUzt4lx2scfbzZxiVfXaCA6s2/q4CsRJDJPrfGkc6ALgHBMRHp/Uco
sI0WPVJtNIGplCunjMxcPtwe1SLzWk3aOc/Orq/h5CeahAF8O3gOJB72QE1l8ZCQYRwQjXZs+2kP
m0Y38A7WeJmGpykHa6ZNmp3ysz8r+l2i6RBdD9krrAwkXeuwvHE16O2kBSfn6zDjYDYhSZHGHsAJ
OFQz0ZciOQxYePDApVGSPLUMwI8gnaHLQPLYvpBDDHjfiE7IDF8vISE7PSxIfurb9n721iDf1VBY
EcSqUSK3f0wfEw+hvosvzJsykXa1V3tfw9rS/r8QTeWPyaAcuS3rT6XuikDArfjlXmBjcXow2PFc
ZRmXHZrZmGE0LvZjAU475usvhRNzXePA4OzsCHxLrw6qMyIe72yTT5nmJSNhwQsBMdrQ7sCWhHJP
87Ei/vtvE4OPWqLNOpwJw2oLikPZza4XUlyqdDutHoskH7IUHv2s6vHB1NYNmdofoThE50hKzorV
4yqD8z+2OZ38LGLfQl/mkWAzOA+FYMq8RGEaV96FsmwFK72Loi3e4ec5QAjF/F3HoXaxxj9wn6ts
fDOyyfMe4AZW78YAwovQcu6geVklfMonglg0oYPtNvzuFAemveNqq8LZK5k5oI240ZOCF6Oa8sR/
UQZUb4Pv+yJKSrk1QRu2qtnhFmIOOUlSf7Iq9C8GpjPjpPBFHemReKgEvUMHPvRZh4AXUPjkFNdf
6TrNZBonJ7t2vT0cTFY6JnF8CJRqt3ROlY+15WZOMzupveNGlPMt5UiLj2tyF0z/34hHYeGN9CaC
Iq+vgk6oLnYfUYlhxzHfz8Bbjpwn2I5ww6Po/k/qnHMdUlCa4r0KZ6v8t8JA1sWa1V8cxy6X/xlw
VFhFXwUoo6rO9HAUN1CBGoHNNbcO2WcIABocLPXHamalww1HmILfqQuCjM8KhRSbVVoXWKDrGmaB
h2UK/seCs+dxSGaTa4sJRi4D/z2nWtCu4D/pOiCy+A/YI15ofwJdOe3pOPpi7j7sEAgQRK4+Bz+M
+EQeONqHf8SdxBJu5BymOF3qOGIb5I6WvFmZEa7I8kt+TXzN8f7ee69HnsDrdaF8oHB+D7mQcN3U
B8CkSGtpt8ELgsPX7YUwMKJ7Y1oPUpuLcJTyuFcI6IIdBE98PazfJo0wy9juMacvL8lw2OrdigwC
kFbsC/ayOCEh4Nh5Zp2bOB96uui1L4Tl4pIDnoBcszI4/EF6cce/QtiiAgtA0tSzi3YbRtOT1cE8
5CPcbXEsjnLc6bVOybzzZZk39GLAl1b6DInETPz4p0fYszF1N6TwgigOqC8X+SPlqXV81QwdxQ1k
qIl7yobw/S53/FeX7Ah55NtsKq9jeXOxQYd3YMEEtaJbwSVkSp0ijeS7iC/qddVjyG4fUnq7Ruh/
QCpaiBlhTliT2FE16B6BpxlIVspnFifropKb2TsZAfbyeO4hYs3mTehKom+AS3r2dtaaNKEr5UV1
Ks8UsnIBmtFWYW3IGOs+m2g/nXY8PUxZosSDAzWFdI6nXzw+hLWV3JqpGljMf28HG7IKcCs3R7r8
LsaKnlgFGYYiAWI7RsI0HhI1MVGxp4F/Z+y7irpRidSIwUbUac/Qowjixr3eWOna6oHopDnYr14t
oWnHSErgOhj41Vj5UctDg4b/qYjSp9+in9q6L2jYTF6d6/lecVksCP1xImgqmGjNkTNHMiCzkugq
XOtJof6JfjVPXjbW7QQfJpF3v3ub1hEUyz7qZWI8bf6W14qUF7K4zeNcs+nDIqo/UB/Xil5lqJyt
Lia82Vj/E7lB7OYZj+pZEbp6xRgFbpaHuNEnel2JM3kfgkwgOboBd/csQIUOPogj5yrWTYqSQpZA
o790EsKZj7fRNa3lY3mOvOLoGTS6fu559pzTrr+9+O2nSiEX7aZhqQMLA5MiEhA+JIX5aZTnng8S
iFs+sLpxuUzkEwUXdOBdjIMwUKd1iP1xXPKNfvMk/hI5evluR6cZUJDPPLM28CnrPyDH+zEoci6m
ICFMBpS0QhqzN9agPJIECl3UOLK1nGJBjAlbcgXoKPLHTaYnFPWNAUyEzcfKngxfKpDL5oYg9bXh
9WVpy5+0vVSn8G6gvSxcxVOlYMSSqcfsByKLtQuuJ2aP6y6XNpTrVSYIINz6BHey0VJAF0tasqOA
IdsOe8xYLO/GdgSHKwJX+Z2BCaHtkN+76RcOosdsbsHczwXxTbfD0gwVus1n37gZ60+PWMQqmyTo
8Qmw0K9umWYIiwcwAL3WUfF6XkpWkUkx2d30w7iX5VD/Y7pUEJb03O36cdT/SK+gYgKaeVWdgy8B
LDe25Hr5IOUltf5vgN+6fKhMtvTVCMnQTU0A+7HwNGNuMfrFY0ZakgbuV2Na5UCNB4kgjL6gxPrA
R5aR6OmkgDsTiac/t+2VftyKfHIdzTEjHpP7AL2jhgWnqFM0tQx0HjRv8+cz2x0Etoh9TbXH5zD9
cL/v74dVsBIRiebM4j8ejGcygGRS4nWoXeN1/Tskk0vJrBSgTyQ6pEHCAH+67kn/E5IqGfIDXxk9
msoKyw/DhTP9gbKA2piCIUVuLV0/0YNZoyB1N0ejgb0QZ8nnrJFjp9PBRdYp6CbaPQewsTg+ckN+
uk6/OtofGL2O16CXL/jOo438dxdlHJYg6k4zBpNjn5WC/VEPq/e9WQJUtclwRZOn9TwZWGuzRPZD
SKIgSZQFpGyX9cH4YsA0PUBTEeK++HjNTOA3BicUf/ToH9BQNHpwFYtYLm99eLzHt27EKIWn9N/C
W7V1fTa4B+gOI/VTDNGRBEnuKeEhSv4cImfMUzkW5gB/tvamb4IgI/AbZB/6jM4t3sgu9VyFp6Ns
bE3oazUOAvJBSzzsC+m0uWa26qQglWxbQHD0F/UjluaDswy3i1tka1xxf6ZzbZZrGluFwLUqkthD
Vnr3wOZw38B/LMUSa6sG/DnikWOyHUodDw19SZQ6Sf+VkPHgR6HMMGES1KSvKwYqRpCZujCRHPr0
l5HiiEYuNardbq6CpYWOYKmr9Si2Tx8tam2XUjVyxr/ZXcVhSJmwWT/Qs8jdUJZhefjx+JYkI1go
QOoHxqS4+Rg3TD3nXDx7hCaDMLG1I1F594teYRHhNzS1Rn1MY/KThG4E1n+nfyn+4nY1qM74/mBQ
UMaSo64n2+65oC89xWfW02XDnSQRcmjF4xoBTUKpJVRWrSB5hyId/Sy8xxGtxWj6CiVXlkOUZDqm
pGzDgFJv4wj8xHxS4FlVDnpSizoBRJvclyU4Iqn/BRcGo1M55SqBMeJD2UFWAHwMC2XhS5J2VQ0J
4wHlpCXMv4nK3sD6eydMErhzkEwnTZvYJXAiytW2W85yj5fNv6ziy6L99J9bL7Pnm098RsdIfvFj
09CWmNTiJEsG20GvCkVh+xHIxNzgByIeN2QtkVDVE90nElk7cK38/rXaPA78KEAS0NV+JOdMpa2x
f7OxceXDqXrGhj7Kop7gwnpinJDM8ZR9TNI/V5wYsxKWcZJ2wErMDXhICdAYpj1l/3wyuRcPVFMv
pitDjZ062EmecVD+BDoBjDJ+H95mb0A8mTgOHlEfyNz9f/Yn8VxQkgdZz4XT90xgJfZsoxqj1Lu5
Gw2d1B5RewsIANkdMivm+9DvY8JCt/B8TRjPNjT+ZuERXkfToRSmDWrnYZa8UwIUOrAxahiz+OyA
ZLnnDXS8y/hIL1vgmP82WxlFdoDu3VIxgev6lLUiwjU2e+wwr2JMeG/zOcvHTrCHuu1w4sGnFNaD
GKGnn7qJC3PncIG+BEWYaVHG1QRTPXpeEzTRncb1TS47LObGnIrdvSfJTbKzmBGt0csQsIDv0wtu
DK9QOvXmIdIfhxhUZe+yoFmj2PGiIJNiqZNP46Jr1Fa/SiW2ogG1/KM76CyosiIWOGMUBNET06S/
VHY64ixwrSzHwh9O0mGFuij+ULmuM57zzq6Posqwxjh0gFNZPHMq2J4HmjVn50RyZMOZJr5WymFv
TU6tEy8K2wDbvqT+ayKcCrSbkwlC7dNZNb9Uvo9GWSdKcIq9eZO8Ug3TzeuNtTThRlbYlUbKLyoh
dLS7EXe4OsKBD3VNrJ5sOo2eUHxQIeviG2Yb3QZMOiSDQj6hQz6/KFmClzCwlI2I9txeZcR8jWSZ
26YMC/B5B0whRBF8X8NXYbQUyGPaK2G/4kgEGCQB/jwWz83gLsnAkw9wgn97oWjJONz3krbLeAwo
Ci4xZen6pZdltdatgFB085D/JbQRCfe2jc+hKj51FbuvDsEkYEbr67uvlWr4vnGFTfZ9KDIeY8BS
/EpS0K9HQpI2KKpvHlTn6Qn324x/xMnoEikvUa244v5QhjXjEEzSyfKJ5cfSY8Wd75yPJe557vVn
BhA6f1t1a2B1ZJqFpGcSnPdIM0KWYBziJgigPp0s3DUo0XFKSarK3FyqGNNjc8RpqKR8NT3FJu02
/jQ3ofEXiA5+/37LbIEPUpYm7cfMdJz17zwwR/Zlf+nv+nL1BhzaP2D67fpZbMqz4E/AmmRCpQ1d
FJvy2joKDyzT4xIDg6Z3oEW8UWY5wsNhzt04N8khI9wiRUsCvDJOpL7/sEwdMlxvTbixUIK2w9Lo
hDQvD4uuafHiPcdx26rsIpy7dvSDmU5z0Kf8zW9rSvWmUD9YkOHNwtltA3eKJ/T0gkfM3ftS4qM7
xcTT5SF2HPuxQIxV3kox5EqMYbsz3nwvZr4PYIPHJ1i3ViwbuhylQ3sgKjYSwmshMCuLCdSAJ/2U
XkcEYPI6CY7It3LXQCTkur27C/Dw+FVg679pLfaeNYhakocuu6lVHVfbMRA3tQ7SYdVmWIgWAli9
s1U21F+aXbHM8J3/W4273wGxyKCbHGFeBIzlUdSKDaAuZLoEjf+D1+x8MmGMqdUuIkUvPs9ddQdH
+26NRvjI1vgs+qqLmO81yIwGKy57RHKsN+ftMi+IwhT5JWqOJmJxHwC7vGcO16YXG+oR9c2fc8Xv
9CIhLeLnHiwDjqQutVRZKHB+wsCBXU/TBvQGLIBT80bAw3HfPWbMVQKQXvVPbuKvvq+V0EOJRkV/
ZoWzyBNhxfRS48oi+YhslbarOjx7izEWiTrChNsORQ6Gao9o/ghBNbppkEHe3fPZusahHkkUF5s2
cVOIabj/HIjGmRAgZa5FR4a0mqCkGL1chX2nhNZxXvvFSaPm3pEMIrhWNEWF2dCSSr4zR7G4j9qB
uzslZSOb/6H7FCvZSA53CGfDCEOhpeytVjlRpKTImZSAbMVUm2sQ0n85+VzUhc3rkXDFqUC9ruMD
NYpNFix6QFhP9x4fyXQpA4H/0pNTRiyAg3Ac9pxTJTwByiYFRyLJ2Yrwuk+ekz6xFbKP+ldDa+YH
j/CzCoQVbVaGGkuX25BUl2n6xs7/oQ8gYKwuKV9e98hm7zpCRXDD1+w8pOa0PCpgjOdZJ2f3UU3C
II/qsI3zvO5r+Js4PSQLVbRPxCDeV67nEzV/m5qUvAs5/iMKYGTpopKVPIpUyO/XSF6WoN/3zMMa
oNdDq7rmLfBBURgwGccj7DKzswSrRwHhrJrlPfexYGfAb9cGpi2IpAxspNnBabaw6pp/gObNbiSq
j6mf6isI33J6ULPN/0geKBpVDIKZIA6rFDgLkXgsG6i/9p04Efh/3XsrHi/4Yw3ycf7+7cDL30yG
ws6BH6EvVGx7jTrqGwomE7AjEJG9kXXW5IYV2H5y+WT51ODiDGMF15WfXKarE/8nbezuMYp99HZK
jkEcHoNz7pWltE3m53WcpquKSScaSKHigzoDNSnfhv5v8fo67QLUsWwe+SYeQV4aHjckYThSgdkw
VV9KKJEk8Kyd3Ae9BE0itmj4JcopULhfA8WZlFrvuwBU3OE7CJpLGSdWdx/8yOeb0/kE5WyAiDTK
B2BGR2Xyn67oKZyXyNN8RAJhtVxq9VN6Q0gussp8s3D3Wvpf7fjCasv9NRttYD+AuSN10fRRhvuQ
H69yBhbhCcJrlfMdr/v58vQWuSw36aGwpfGfOFzqQdzfJTXI85UiIGwvO9Y9G141vTcYXCcxzH9M
N/h7dykmdh1KakqqsL3VKdDQo2Yzrw7rcjzFD3MvazsdyyxnL/QQSi2XQEdDCyMoHWht2MzPRcgt
Q6Kx/L3m1R3ychCs8H+J9CfboyEOtf1N13QwRORzL0xoxUcd1noOOjGuWTgDyWDeoe+oDVCNIk46
TXXQfMmaP34UFwt78fhcpaKB341GTux+5msQ3UW3hZdz/YQh+gXx4h8iVbtg1RWlfgyodcwpHjnd
WeViqpMOJRVHxzEWgW6HhFWUswGLqnD21H/VmboozN5kcg/POlO1VqWBXaGuMeuB5qnKtOzyoLZZ
2yoRZzsrxl/ohI0dt57nKjVCweXbFNNrHr83hxZLot6//qi+ikuhxdqyu2geAc0rNbGSS9le+nuK
dyv3TGi3etKNCjCrQFAeyayEL4KAThHgm1JM/2b/8vnTyPERuYAWRbf/aIj5RP/JCn3cxUBF7Rt7
XfP0TmdAy5c7pInF2/utm/ZddVQWplbyeI6V8uOhkBpkZ1p5DsT93DD51rrsmEivCA5MCg2Cwxqp
ZHVV6zPogmIzSno6vKSo1CbXFTUahexRN7bvWAwbjAxlHwjye7vmb1mO5As3v0BbtPE4MP+6qhnP
DQduj2QCK4pzpnNCOPk3UjpRcagMegOO9T4jmL6XMkk8NItZSae9URT7EUsFEc9FWCTeZbPVNyz/
BKWbXVaRoOLh5OxoNhFaasTTn5MZDEJ/aSDzg8yOYNmps5u+tE/YcdABSM78fyMvr+wF8WsqodVi
wrxBvhc0+MgRSJ6ZW9ose1STr8S8ctTnzlLz/Ff5hqKJ/HL5VdNlK2NXyZg8tylnbXJsr7kecwSj
D4NPSZhEVZju3jnb8CNrQjRlYWQ3oLe1WstosauWEW9tQPMG1ak/d49LENJsTfPzOtXko2Gdxt67
w/cTIC009XBWdoYAC81cX1GMqHPDo/C/Ga5uUfQ4bteU1qRfX+Plw8MvLSp/AQ8/Mh1s8tAxH392
IfaFtJrsleFBdMo8w209bR1180RLlUTvNarpsMyvWg/01AtndprLeMZ4pNcOATKuQje5DzVHjKEQ
rYxnRzv2U71U96oRcuPJBo+Kf1EomRmbL6VIDtddkW+2jZaFv0GhsvJ64Zw4R4+B/MqsVBc4cbCT
6iGamv9kp3VuBshV9r4dNrrrS+qAUdfoV5V0HB2dBJMs7Upt+opAUWfH9MWJ2SH+aqtIaYbuz8Uz
BQHc8LwZiC1vDKnhNyWAE9HHb6LfXhPV7/1QP5ujIY6Esg2SigQxKZAJA7uleH1htf/Zv3W/H3Gt
j+otsdp96Xx7BGidus/+C9VDO+mCgPrD20lDz6SGqBnTtLzjNLxmxf7WSHdJRvqJIa6KuesbcBZ6
WPuvbrCJSvXCR+KkHFoYo1HqoSvSsC+0ks4H5EGNQnbJyH1n7iXJ4R3XefIqCKp64FJOuxELQmjH
hxOkgU0WxmGgu8vaI4WEFIOm4ORmO7AEQ8OD/5SCpoGpu9utNvBUZFGNnIg5cB/mnITedL5FSWtB
dfbxpPlJJFLgsn39lS0b02wI7DkOy1MTHNjnIydw91Vo87hroEF6wYnBVAihqkNqsFaCxByGoLUi
C4MyZC1uUZZlHaRB6+ckZdRYGhuptbf8BaopDeHlSWaGWU9yudrZVyRtis1t0xvwY+Zh9AGiheEE
acXepe06fXrZ16ttYTIXLLmFl0du9oKkxQk1z7MYXch7GCYtKnrJYofESAr+zKvVbltxGq6i279p
KBSGTo3IsSahUi0tMRPPcetLv9S1t0XWcxiwUFLeOEBB66e+VnpAsDsuWpVs9w6pNsndnnYONrJa
92x4AmOelZVC/2PpeNFqvyl90lOoEpeghKfSBF1CBnE4HMGnQGyTCLTbGCmLvKUgar7cX933/SIs
wm8BU1WUXAiX0rBKpq0nQTqMH9M14CKvN8Q7Q5aU4XQ/tY5x+awynudZyQ60sVcAMNHQAmul3HJi
5GVxizgyd9DI/xVlgQZmryGrBwjDLM+W1eQUWxGDXOuZWYhLEHXD3DMyYWeLX4voeBXEcmV4jYe3
PVXh4TUzggLU8RalSrEOp0bhyX73LuPL8AI9kYo+VQyqWYA+8SKZE1hc96eAT6lwMsXP/xlk2MVm
XdL3N3Y46x5bMdzkVKOhwDQ/YA+Fsi1utymPpE68eTWjOIVpy0S6SeKZJp2jSTzCu6XiRjRVYXVi
vL0Z0j56dfhijxoZ6JDoVS7Eu8i7GflC+Y02Z9AVylNiWq4oLocJEYS2Plia8d54lK0CFBjOgIOQ
5q/JTeWUsFPjtitkmSfpx2esOc7xKFhlZ+IyftCG2JNyXXViLl+CvrDhtF+25hky8cVqkV17KaWX
wqFS2LqKpb8RYMsAZn0+WL1f7qPv7wiZxYKfqXtmGsR//mBtWS1xp0wN8U7ksBpAAN8m98Z4JIPO
YHSChbYYRv0lpt2qCyLnfx/1OuOEbHC2MUcvdmZqzxpe/miDnxNXZMhe/bO8etd7MeKRD0TlOSPe
3egKNY9HGA1CItlGTshJVihcbs5t/Jur/1Z4bZ0k8pbQnM1ooI3kKDG7vrLI+Wb6gieUkpy6Cjee
vMrqBACxxiTXE9wEanh7v468j81SDQPheaNPmCpDf4NDNL8xM5OyJV5ZvNZYy5oZtsDkSjSl0v+w
y6pgfHhvWNkVsDnqZcNwKtpDEdHSzNy16Yj59mJX90GZRC4vsH7MiDqAiE97+1wvqjA+oqGdLdc3
Jwei+HzHMI96N01mER+AKaMxuO/Up2etAelrba+SOAxTbAhMbaHzsznIufuTZFi7kwCMApsK9MNq
M+ucRgfIQljajqxiSnSQblDfkR2hnVRemSl+XK/JT/fdXSa+9bvbrgUmlVd4AapZ3PWA9OvupK21
yxtd52R+xmItMizT4lgWSEXtNvRtzTtrFMpkU30ZJc/DpeWreUcRdhVfoPCFLZkHah/izrVgYyoq
Tc4Az516GmnQv4yC4ZIUi5r8E49O75GL5W68yaAdmYtsi6ElApcL7vpRcRj7dTRn4Omg3o0E45No
gtMWcVlSE/szL7qObXZUA5iYVNWoHM3PbcbI8W4ItSfdu4YoimyTXMmzU6JfbgU/cNkCnpdomyW8
wZjCSFpJFcl4S1cD9yLr1nqGhJIewdTSHo91Vyn6iFA4tdLsQxUS3D9qyb0J3L0B676kc9BokZlf
fH0GGjOTbl8IXaMBZ3LeaRfydUvtAQEx0WJrCy6PcCP1EdZCgU/co+dhtqkpOEmtVtU2SzTgQaVi
IXg8RLamKeNPcIKS/b/qJBoMkIZ0lQ+TSjn1jZUO3vTNFPHDcT+qBZS2y/br57ncLo8Jab8vft0e
oSxaslBGcsm0NA5kwE5WVxrMDLdYXgcfsOWEa6Ysf10pEkAyeiAWjXtlI1jjw6KE5XxX2dyLWYnP
d8uxZ//b8+LsvOSMz3IT1xRaMB/9YIagqxkommrYppyF0/B5GwyYZc7fcQiYdYKeHKMpzkkbqP0/
lPJuFVyTXKkf48YsDOpWjd6/eASY7HWnc68FALUdd25Din0EOqLZRWNFFuoJAB7LHGHd702MgkUR
k5GXWdLsxiGTEQBhJLhIGVwQyU7Smw61PdRLHxqMDStqhx6AeVoDIb3BYm6mFNlDMFLhLRf5UIxd
e9LoXfMokY30zJrVXlKVvC9sqv2MXDWhV9SssQlXXYqLIfHGQev10QiE/35pUKMk2eJoY5HY3Gkd
1hARjH/4HCjGKJu2w5wtaimnyOMT5ih4yJ9LI27oP73ASG3YTgL4csP9O5LuCYGg25HvC6jpcJLc
vrsbEQnfRXTcJKsffjoUaalt/wtoB3y3szc7u7Mqd+1fm+/v7p+Hxn8D3ELoYKawnHZtaLXGUWCo
jT9SBIkwj5PP3ZcS7fd4Kcp4CbZ1PMx81/p1Pe71BZ95tY1oig5yh7nUn4XM30gjWmE3USoW9cj8
axsv4fPx5rInEhq+JuOF92+NuwQtmcgzjNSJsdpoRiXtVOjzu/wjGywKjn0Ssc25PUiYjDJN9Z/F
n7SNI646POylnk+7I63juROuuH9eD0KaOiIrLaR4VcoxTDsF52s2oHBdaAkx/TSkhnW1TcYIwcDr
fcj/vdn6aQMYaY4MLeSrQzbZRLbRjoBH+ky3qV8O6/QU3v3xv1t4UyVHmphzbhPIqEFca+KbCzTj
GgxOr2F0h13/7k7YkdSWojYkBj+CKCRNjWMjO8TU2NpnbMSEOMrCXbGETnVghPTzFp7kbsijU6zo
+lfIgfElnVvYXxp2/BOY+U3lVx+IWW89LGGF8FDLT6IXNNFpkWCaJIcMRLgn0SSb3OwmbisfFJOW
XBCydQvVvjCRD7MXhvxfjLQAuTZmlt7A8di8/3sDpR2TduuMAGbbx0lvgByEMFszWc9uV7VgtQKe
dKT8jhw05jBoB7TW7l53KL6gh7baxIsMyKmGF6fXup1D2DvTo38p+CJ6glcJmfTZBWuH8MK3s7+9
GItES/EgsN9FYDVmPmywccE5y9pAk2YYSqY1ot232+Eks+yzZ6aGz4GbaeArxhPhoksNgjFLz0LU
qy2qYgDLQMBs+QoYtfW4ESjlgUCmvAC3kQstYm5szUbtT4KF3CNtusuH1olyXFqGWirefP1zzSeR
03uM+skTtC5ArhVWCOozG2w8VOw5p+esA40h/WTSNVeHsAUvHWPgI9OsyN2ScA6ySdR//oaUmDD6
wBajrXyfabkbTc8VFjfjV2+6NriCnljtkWOxifGcAi+1YA+vMleElUdt4icGMn35XGU95wzm6zNR
Cl2iaAte+Q8p6Uzrf+lVL4zEAjkBupdZqpcVpLVJI5CIjt68RldLkvyHEMZT1xWq3TSXix3qTBGC
E823Rzl0V8M4XAfA5Cms+63/Bu0eGBJtNUAGPGma/NuR/9tBikSYKECJImE3Z9TrO4AT/jCUO+1H
KOSBti9XY3iz16BGpJGjhHaXmQ0YiYjv+2lKqWEPBFR20ce7cKHpAKMA+Q06shUQVkJY7jc4588A
+fqyGf5xLgEha3fE2dQFwfzbBTqvsI/efgFohppR+V3/aN35eFP2aahCscVNjWe8lv9Elpey7fjf
C3vhYbaMqubH8h8pSbD0OqfZncxNBLzFoldfS2Tg7tFD5Aaac5HEForUciYLdTeGs+LEXMt5yYYv
qGtY4Kks14LNpm1Z8GU3Ux5g5BXU2riRgncsfcI5c0YykgJ0IF9nf8rXMWi4Cc4yQmJfRyFi4/hz
zHR6S04PFvriDEexJq26ut3nnxQRTwZGSwWJ1VyBrqA1PFZZXWtaP4xrb6wqR5rPxycTDth48Ouo
YwcB+9zXBSfg9cnryHygUrr6Kc9lTcxCjAeOvsNX2WCsV6b8MLnVpyBW8llFqeo9v2wlL32xObq+
KuVY1seBOOjBIazXw37a0nAiMz0zodx4SNGtLaRcXzVQ2tDneo5IiE6N4bGdCRi0EtXlpUE4AKJ6
BEddsi2Li9jrpzkn3fe/QOyBQqY4dSOLd/C9x+aIepW9R0xPujwVtUnjk3popM16zBXKIhKuIkzu
TI1gMtxYfPwOfU9xSFYVBjeoVjddAs3VL6mKP9/DjNSZXTp3msOAAfjvEZLjhjxfJX0Fe5Myy0T9
/NfP0l4TYECnZlyIKbSrzWk1E6rdD2g8ygJsvg2nV5WeiOaSpFGOBqm7tjj6OlLqDymcMDRvl4J2
aTbfImirZEAmU/t0+GKx7nb77amBolh8vux38ykBvxuyiN8g/MGmFboNdOb3p8MsXXOkjDLAM+xO
kZb6tHWPxB39ILEn1e4jbT+XciuMoGlARbSpswaM3hk6A8MlDLzY4aWcJU5+J5ztFLI/v0Edbs0r
maQPBofm8Cy3xDBnCWuT3zjHteNpOjAL+PiLth07hLeYT825Z0hbRI+btRMtM1uGcx2vGshe0JDU
Fq9XP7GcD8jq3SzG7mNM5yShC1cOwxOPhaGjaenwFVEeI5KevFFPstXaepaH8PEBIKsh1mI7J20a
OWUEscTnwuHOaMzYvF+Mk2akJPCmVFX2T9ZtFGPX41EVNoL3EvVRft9GyMVkS4uvDFN0nuvwrcjy
1PGBKerJTAH2MVH5EIAsMiBl9znkCb9wasDRe5kEU1VPthQcrOXpivNJNfQ8morLoQIjkmIVppXV
mE7AqUVbrnuPWsoS91UJSL4txvxFilE7vpV0ohAEZYvLU83rIEd04yDVWORHjDYJmSAjx7p07fpd
53Q5uLXdm6mpGIPHBiD9JPFPFTRZCXNwFMbZzMBoNz2LjmDfFgamomzwirl5/dOtZATB/TX9Tf6z
SRdwWU4lQ7pT/ujLlS8pG/0NfX3A1cLyj6VEL7p7UMSpFQqGsUMRBKI9+cmtKWEjjVyTgPBjm4Vp
GepcNTronfln4/H8Zw0cHTFyLficHKtcujtcxsIkbnt5ZUn5L08Yfm8tXrFpI1FKhBriMZZHKJov
yvm8pMLeTUZMYwEmfzyu5oqajerPg+18IKmaBYP8i+MdW/xyAp9db0aOM7GLdmII36SBXpsvVRKS
aTHVt7pp5HBPkIdh99wC9bSs0W7iAv7aj5fDMLWmnwAm/rnSwdEz1NxYUkKhtOt/HDnzKoob70EY
48RhSS1UtxSxw0ATNgtvgr83m/egKi13cW9ddar9pAsnOsIW6FkXHLaNcSpyfQm1X7uIaWTkAq1D
qeuyYtnoGnhmF5lvn5VmR1P5D9tE9I7UGiIAXN7vCFIGhyT6gFRYwZyXQKcSldm2QuEbRfSMqrAE
po8iiV64GkMTND1HsNYYSS2a8uNPMp5vQQQTc+GSko9yfRGFOKloPS01rofMSFmbe3QX/Rz002MT
lrNZtVRyoUelbbPaQBkbC9Gtjt7oWXgg9NvaRPs4PFOcC5RNcjJk2mQYkDaOogulmtPLJdbheOsg
xEXkPoilaxBnH9BM9th0OyooRjjVITsJkHn78EdO54ZMYpCfm2bt9YTNncroUPW+H8WhjWIAxYLA
LASHcDMWptuMhRwXhOmx11cBOkFzFqAC8MJwp2fSRywL4gqawjHSmFxVbJikNZtQE/8hwgdT8Pgz
uaOZ8yez2aimWefqav9ocBVUTnM1ylZrg/vbNmQgWeDUkBxlnP/t14818M0NErDqngH7zNz1kxp1
YCFQLggHBzziLshp/6iU4fCEjF44EzeRdtlfb3+rj1NyLbjYa9OHIZlcb/DYYjgMtfHtatEa6cF/
Nc4z+jaSEGupN0hHmX6Lo6lHCsmwtD9k+CZu6fKBvTnpAkmgGa9LZ1Cxb9vyI30zKF6MAerlo/02
V+QwdAa26KzN5Vu6KME5H0Ck6Uw7ru0W//JsdLvqiKvR2U1xdt4tm2HcbzWYCojztcy/NqfJpZaf
HN9dSIfkHF8mAUBeD2CQxROl5ju6KMptd/2ypctXv1IFpAHjG1QUBKsw64XGAkK72fhm8lEaQicX
smpGDKK1GU7jj6rFbNQN9HE0Ed0Qjd82bf0fiw+6DVJis/6YSbRELJjV3/EohFt2+55WfQJ+hFz/
Iq/FhoIBA6r6xGI5nTYuLmP3cNIOHZEe0AwflNoSFcbRqbQKgBVclfWFFPu1gfwD9bxZg+u0Y2gc
0zhWvUcEaT0ATY1nrq+FNo/aFYILDd0f6DZc4vs/4mLn/dnySVOQMSkpTTCKW57nTFWfEPn2FJmY
eYuO9kdSO0xID15/jQYAYR0Rt3nIBxjKw6M7FjWSHxNKJIhLBGtNTTJMOCgWgvtcy5UWBsWCNCfh
ITlhjLIsUOpgRU4ArahWhaoKdajAb4lSmGHnCPADektTD8JDYoKeyqmQyt+L4/CcrAbqndu0yvGx
tHsrO3UhEOoZ299PIINmaiqFJ18cd7QS8IUgh4gqiepsMkr+nrfd0WiuRjveEOiFrh75sBVgWgki
6HO6+iNbgQAKzaTaqrSw0ALUgeaVG6auXGOAXbyFiSNPNjj75O+hyym6CD0KtnnSyEaogLbVaL0Z
SYKS18p2A2Z0azTUIoHGfq81BKPvtE/q/2KY0lDf2WwCgTrtCuU8bF+hZjNC4XFdhYNMpHJ9zba2
1a45bPxu/fEfnRVc7f0tKh4K6etuHvp18hF+yx1HIbkkDaSoiv172SH4Ct7laEexdddS6Fz7FiQL
BzgO2++qgcqa/EZsvrh2l9EV3U3YWNmFm6Z0YBKAWIEZFdDV4oSSzBvxr7N+coUwAjOjLRiaQW0e
KfTe26TJbWqRMgdVZRmgBdBoW8QDtzGd9IYMoub5mijLHc20yh8QE5MVrH3ZatS4c1xXZK1GsOY7
Bpd4YibrRu6ajkFfpr//81tL4/RgZPnT5TfcU9SaKyO0eZR+8MaSbfHL8U3knrzn2R3ur8LIANZI
wTS10pd7ydUnx7giRm7qo/aMPbSTamTZLT5Km5QD533Du8+CbSrMUE4hbCrS2zRNPP1g2d/Jmhkw
BHtg5izFCJ+1e2X6k/unISNj/pvfIqczLBNTfSd1QrqaImT+2HRfuWPSaoBUpmkig4k7vyj0cSHV
9NcJesqr7XoILVu6y74adBw2nLVY4KcTmf+CFl8SKrinpzWqZZgnfNGUtOc9mH5tTB4zvvxprCJW
w4A7O3LGnBfOcdpDdJMadZ6duQkU18+npCuKqHBD0qyskRw/Hysu+ZvtiAU7XzRNEK1az7OZKFmQ
Zn0Fsawma7Gc+X0nmTnDuRuXjHctO1ZYQs5fAAcM6hXXwR0JQ2OoqWTdwkf9f3DuD+gus3gcd8Cn
a5OKc0Wrz1Z4CLrNbtC6AgRjukomveK/jEiqYFbF+6dQy66FfIFP41xia0iAyMymy5bckaePvpFx
vdVxI6npDAmGzlcunZ5MSDxp7Mqbc3igCFHD1tMIJPA4DG/B3dGqI/4jgxZCkQu7alGtld2FYtCS
0zypu7euElec8MpItpoerhyylCROkiA70e6j3PJF+Pdn+pY0J6NAg4/5jvf+i11VNdKBAXH0XOi7
K0GVFyTzNub16KAqdAYxo2M2n2G/FoUG0m8LcIUaXhHXXnYTEnmJ9ymUp50M6F6kV4a0L2ln34LY
YgyA19Nr/cPMOihRBPM54Smkl3PFA0/oC64RwhsSKVPgC/Fik2/XDMNUClSV1jm8GDwx7MP41ywc
axtuDtn/mWoiHEK7LnkUK3kizK/46FHKoGr/TCThpdPPBd5lC01dgCUxVEZ2u7mniQNeIAgb4no5
+xCnNiuEqj9SPhwe/0ZM/J/sViupjZYrAIU+NQ/DHme1WsOBCffo7qQcPPc6+Hosrw3ffJ6Dq+Af
MsNnzt2Y/1sr8GGgmt/qxU7qYKv/YdQ8VjucA2FW9X+/+c83zn5kiS9Gdn7y2DKYrENwOfUXxSmv
cS3nr8ThOYTrG06BhASOJGO6Ew/7biyYy9s7LQu6gZYyjxFH1FTfQdeb1nsGD0kVSG8kekcNVHLF
P/wU6SysN7CyFhfbB7HCERtADT68QOU5z3y1V9yj+lTfa9LeXCI3D35A1Z9E1JJOfk/wj0h7BH6o
KTmic87Jl27x2pxz+hmOIqtLqUVQHfnJ4pHwIsEv6A7J0sujXRhl2uYP3HGIdYrjy+yvodYxszkf
SL4wqoiCBYneJNog5GIBQgzdtdJ/KajW4fyOew2VFll9kD7608633FavoqMiuYBFnLXN7JAOwKUE
LNe+ld6tEves6n81cd6kVXX6aDqtiLVJ5LHGIPSrTQANg3ygkdXh3SV021ZuIaw/1ZyjtlO+U0EQ
+8w4dN8FQoDExmXfBXecObMgxfXbty7jq6qnqAZ809Yzvh7awjfhvbTLxzb3o+nOQPg0sOF4Tnt/
d0TpwP9q86M6ODNuS1nM5zjnDMGfsRg5mI8FO6qW62Vs757uVejGOYZb7UYr4nM3GlimLHjxaLy8
qZfI4MS1V/U3t7yvNKW3EldTAcmBEi1VGo4Q4RZhvY57/PAqDPJDPjccmELxtVGGMF9M+jjHEBsk
7IeyAV4WUQsOBWPxjGOUh7EZ5AL6DleavBKZZigI8j8Mp1D3ox895vakl7vTFfybGwlAYfnDxDhi
U/NsR8SgFa4sgJEo5PTk/we/sQrVYe5iqkvXXHsbNRSEH/8D0nkDs328H0+dlSlFM94UggHzCvuv
4MFVk4mM2E4UzlDfP1jTI3r1TPP1vYQKeN502Jtk0CAi0onbTUP47LIBWyum/kHPxm6Uy0p3/P5A
yEt6ovvsak0u5wh3H6H8US/tu6XwHGHpn7TSBfK5OheP0gDUPJ8JMSeRtikzKSYNXlGwd4OCrlH6
dCXRKKzsrDY5pXMXnwHwYOJpRIA4WKRaOf2k44+47aTunDpgPUignoCrH51e2exRvDAgjvRCCctx
+H80wIa/f5KG8n8/r2U3uth40eNwg4qB94QSKWRAcsZJoB5X00/YqDgBvNU/cTS2998y2dOUgPXC
JfhJ6ZYzNvH4+u1QrIHB8/2qBF6YJ8rkG5TevPgfWNK58UXKTgPV4QoLV5D51c+KgrKwWgUDPvio
sSQ9/rKTHS/YqSuvdPH90eN1tcZBB7edy9h/5umghX5tSyrSFvAch47RHE1Ny9fIlulfhm0OSAdN
cCUlmyMplangMnQGFIf8XPnKr0DDEQKk+t8BgLe0w9uDdzbAHOk5TtDJ1tO59xolNBCm4wcIqsU3
y7+a4yQFJMkgpfC3CJ1ZOgKD0f7do21m7GuzFwHwEgjR7O/qhrzIlWIPi4laiwOzNs9rXStxzsju
XxlNF0tZ4btM5L94dcIW1wqU/zVlhi/vQEZbR3Ra/lsV9ytny5kIGr6Aio4JiNKXP9G+7N6zAv1V
CDnQ28q2m0DNSeHtda0IjYBreyF7akaW01pU7CB7VYspAx3rkIKkS2mdIclgNBaHYm2UGYqBAnAh
1IRZOGTMAVvUHGL2y86++3fdb5XWa2YyGypAEpacKGNs21BzC29AbDOFOYFJtoE+9MjX1BiMS0nk
khTQx/7ikqe1bTelNxvqjSW3uwQmgUZCakIZCdifEl/10sAkokpz7vmSLcX8spZS3/vmWBSPo9Ax
eCQGxSN0wy4RxQNbkoQUC8xbQIbtTaYZ1HNjT4A6W+xnEvWW1cs6WG17SWgjNgbR12gI/YqfamgA
HADvDmte2XZwx+Ow31SPTHvh2aTgSv2AQd6s61PjLgClLzva1pJEqz4tUYF3Js2nW9p6qyrh1j12
lsyL+25j2xMh6tBZFK8PEoKFCqAKD8J0Eiral0MHr1vBIsqMDYTL2+NrVa6/y16txIXTUTC6YGUX
kNSCvX5uUDVisx238SrvDlFczOMiiMPTzm2ucfQYB7GbhbMF1vEJOaf5mAiE0Hk0HMJqfWzyv6L1
BCpCUisasb50adVuy6dsC8tzdpQTAM3YbYEd+TllUr/cc3RKtUnYGfDC72bnbbMN+by4TbMdjC2F
G2nxC0O52EEkbUEI284mpE5dt1n58XD9Qkb+RQ1kbqGlPzss68TmI/XrY2PmuqZ543PYtxCB5KY9
ux3FwdkkkM9ZUoPYA2tJ9YPxtH4R3EvrnQ8fEDi0lW2bSbtk+0Kze62I5GK18pBJwdWGYfFTSknx
OQu6YuEQQchOAgXdvY9jSNQ1uROZrbqUBNZ1//jOhzP85bxwRTr4iwi0Dy1DN6ad47UaxfMVQkJj
+4rIHNoFp2q8AVYg3UoPl1DOFZ4dTmOW6nj83LLpkbqDC2mAQ3sLY7PS8+rJynxtodBgke872BbJ
yi34oiYkRwDGmehKCr2egrZoVSWGBfkKhg0/MvxyP7tvqd3kJy1w7nkAw56DAM2IJwEyT5yLoliI
b0t1IX62udeTzTVPydytFFR08Uw/dKlzlhIkcHucLvizg3zmW3o0SFiacwGy5Dydtoz+VFxbATOv
HGLDJU/4LLSFFlFhuB6caSsQetDkgW5I0MItJmfET0HSXj1umO6Cq03bi5OZAdHWVMwev0iwvlYu
Gm+/WCsK4LkcJ26MXCm+PCF0bP0460D//DL70p7G04arGdENlp/K/Ya+IhcfN1eUPlfomWpAtIeS
9sOuNWYJyIJ+A/I5BrkVeFmeqjhLfchIhQw6GXYU28XjZCyRa9DcQc+jOi6uc+0ubJijK8Tp4xSm
0aRTZa/6m1nXuEXZtLQgmKtzXcMjYUl0+CC2IwYzWFUE3g50TsRwNH0Jf0RXUqvwkfDE+R9SZ8ja
mo9lAnQ25QB/60OUbum47qJWw2pin9ZfBQHp0sDjkXd/K8rDKcwW3mldHSYOgjxUOIihVp7B1kD1
+hrOkoM84EbqbXFsk/+8s+APVnU8UrrUzkAnjQ1hxuNYEv9kyGx+jAoThGzW4sK8PfpErkfKdcZW
mRcBIlnioNKzH0owA30g4Y1EKyHL0g6vc6Df9XlIWYnD0Nq/ZwyKexGkCuzF8UFS1jWyplAYZMy1
2HslJL0QGodkI9FDmwNPyd4M7RdbXu0Y5GjyAD18tTo4b4aytEi290khgOQKVBDxtD4XNVl1aDlf
CrKS6s4+P7bwRPclKgmZ6ug/ngYvV+x0HYnbF3az4XkdGEiX8BVw/w7pTWBNnNIOc5EIHMBXQlsg
P3TCYYel9XzSBsvY9UstY4uRfFRMC92XvEFXa1KhBnnccp/22dW8bD+Pg2/vEvrB3IVKXQlQK57l
NGflMBXR0IFrJJVb7K9H3c7FqOHkcYkgWJcktG1zI1zd5VrxgvTakgpHQmtvx1M7w4jR3/irx05c
ovZQHh0HVzYAjFst5K8S3/690Mqk6E/kmB473Rg9E/0tDodW1y5wcD6dMMU2e/VHJsUUwV8O+IGP
FonIBvn6OSQUIKWsUCiSS5pghOWBZcXiWPB0E80W0S13tC0kB+Q/VePoTbOOarGe6vuApe0jEvBU
px96cxwVbchwPSU3qCdBlEzG+7wa1FCj4U/1ljjnD8Qrsa8aBYghAOLQ2Ftah+FGEMFBJqUKkIan
N/qu8sAdR/U/HReglJlPgK/wLbi88t0BujVhqvOJnNld7g+/tgfBWWnvXsYyptBE0Bdwm6f7BX2w
deT6hj/174G462Htxpo6CM7mA/bjvrTAL3fprG/IsEwqb2N8U/gDsY30ZemY1MmisnAgnB2cQEdZ
aEqWbBnUdzHMk6eNFlDZ1+t6xoP6aUQ0qJMWKnVCqnGV/U6Tj3dEGGTsgatTomFMLFdxOMG0988n
eBcj682g6HUZbLsKOmyf+WLiAV9x2iotbH39NM4wetgvtsr5kG/K2iBqSJVMh3b1Surqx5Z+hMxT
x+Uo9JyInT2mcdlb+0TrG97GqxJfinqNP3HqsPgM+48xs8jLdGlu8bQoPKeYm7nXNIseBzvpBXc4
kgMwoJGI+X5My7cgK4zn0OWSbDxXgNV5F1D9H2FNEP9d1Dk5m4p5J35AShQ4gJGuiBbCkVHLSwDz
yetU9xX974A/hls2NvP3sJNMNu/FuHZZvDPVpSH7oQZzvGM8qEPmdmR3629FHp6zzcy7L4pfI+vR
f9YwV2dubghvSWZybtiRZlb9WH3x25QK4nZKwyzGUvubsbn3T4hngWRmQYbqagTMff/++u5gI8Pe
iuWc0OpiRkGHZF2IThn3BnIp2BC7r4Sfj9kb+1ZSIzXkdjxsSG0pbfpLYJZi9Mw/lGWReVR/Mhur
wr43SHJX1nMWt7y2zx6Wsi/SqmKg8HA1HD7qkL9XtUFmITzb3LxscHRDgjuUf2lcqsQL+fJbhIx4
WiM1PRHod7n2jQqlO5G9S+6tI8zJ1E0VMt1/ZfcDTSHN/lhU23+81dt8V/zaAIFxoUqAx5BS//IA
RfnhiWfm3wy65tsJyjeHm26DMABi3a+LTs2byb5rFWiV4vn3zJc7aj0XZRPar5Q1lU9gAmCsLWQX
7dvCGTeDmBPSuy9/fUyD36TDna+3ZClt6X7wVhBFC7c7UAcd5zFg1lnT2AaoDreqtt8++q22j6oc
eDGSynA7dfUj+6VVnaZqvmdXlTTfyYhdeWPX2z2yAkq984TtneqGNmkvxJDzMw0sHb5TnH+6y4Ci
8LmK8rFm08KlyrlbkuSeMExrq25DTEPsaHSGnDGrk+8nxQtuWWOr/VI6mFwFc4HcoUQpfhNqxmvC
qwQ13bWu7MOjS0Y2xkO2/NMgOU52BB6vHF7PDIFlWFCMREPsdW9tJ+SHScyuyNXfi6+e7sMstr9g
CQ+cWUDB96B6R0Uu1FDbOoLLuAszVCdBkSdX4tQ3S2xsWTPIWyowX3tLxymHyPj3sEWcqWOFH7/1
F/iIm+c/WBGMeIg9qmcRQVWUl6PBmzQQOgF4EsyNXig8TztIksQ3uY/jWSyuwdBY29S/z4nrJDVQ
bjfLQMDKhjn2Oqq88GZohe1C4KHc84N+5Y0+jdnJjfVmnSKhtUBAiPFfh8SMzIQrKqwca6xgRVEw
g8KtbkFmw7CEPE2YFkhkNnVyDXsAJFPvbv2Tx6nmuzUHKrUt/GdnQzv169DNX8T6ePXG2r/o9iXm
e5HwEIO0l79oFMvNGgBxA0wXbNcPbUY8TRaCk1ZfpkWvG7SCr5vhQq+z/wZrMoHomrG6N1B64TH1
SyQKZdlcgDHoZzjbs+ngEN8nwOadRtwF9ffD97j1QK9BtqZ2euk8iZD5Uj1rWtaUTSx6JQfDSMSj
9u8lgphymrWfReX4Ni9ncdO4XKNKIGhRMyKKEhWIzTChnnuWi6rNWA2UnzGxuILQf7NnWA03a9H1
ENSijoswRQZ7vHf0erSVNbLXRoUKLkVUn7ubG9zTH6ChjEthVvc188BX6EuGvVA9xbxMwbGEBHyp
66KiSmls4zigVqxpy3Luv+jxei8qhH8/NoHm5WhP6kU788CVrAa/p8Gv/1Ol71YyhvuOo8s4rzax
DHnf6NPqjVvMdH65gPqtNsjzS9plYKTQaDofSjLmEiH6NR5e7UdJ5sWz5BW83zKumXt6RH82R1RJ
rglvJHsue+ShjVQFqy/nglNaeSl4gtLELKF5r0dgh4NzOgu1ChoR2ImTiiIS+0bDZaooraynk7d9
szQ+C6q2trU9S+9oi0Xo+EX7iXryEQZPmGLmzSWMukfRIWJZotL1EqXsuept118/T9sJ++h6QNpS
jHwkn4cfN+EMpNg5n089xX8eXmPzTnDo2rv31eKQqZCDi2+0o9osasgUEjGI5JJjqs/gX5LSGdJS
lCnQO0dK8lJtMZ1N2NqvgnoJZOTHUoi6T7n/1q6reYIm/IXqA+K+l/ZNAv3CmXVHUqrmqCteVLvg
fqmbdSRryqSVGhmomFheJdHNhjcd7QmLu6PtFxqYmkHTmT2zSU84oCqxX+cCwLj+/pv9Rrs8u5UY
Ab9B5fcKRaKlbZczVS3Bx7CTHFblA+iRL1K0Go+hBqu6FP0XxzTTINWRVMx/hCId+JpIoPY+BXsp
I/xasYTfCKva9kLgqmN1tapJsW9Siez+Yv5ZUnRtfUwaNKB27oMRsSJtdx7hGcnYl7aIoF0cLT73
8VA6tGi09x384f8+Efd7WBQsu0QqIcSmfXzV2iTikuNZ2ryJD+MUiYZhcPgm1QStzdUfiCaghg02
gy0oNoQ9sK4amSVvb8uHB6D/Y9+rYgMbnWAablj9DIsMtOc7khJiZvvk3gl+t0HzvNYXDzaLisaZ
aKgiiqXhswMBsSOg271hknaLb2sGTXUDibEtt0xqtY2K3FFj/c/fNbcniabCttDhSN25sttC/qPg
xoYXwRL3C3GxysrmWiW8QTlpw4N4K7FGF0LY9TW5UGIxgggSkxuD0RRD+koVaAN7g5mXR4GXI+vv
QB9srleCnBDHnnbW5uu72lTLfMenZL4MX1+o0cizGBZ0T+yR7flyFfwaS9tho6XWyAKMCRcNMJHj
fygs3fzyNzzPgivmZVn12HTYoq4k7uZRNLw2GODwamMUdFAeeM+dWKQ7677pu9j6fQpleBDEWMKp
TqVNC8AwvMq/1nV1B58w23GfcCNKCih9pPYnM1nULonBsuRK0i0yeLckIjXJRxY+yloUCxK3LV+t
aNSE2hSCuS9LLKXQHgzBS3GuUc07pZC0j/vXFogvtfKR7u0qTHhlD7iBdtwhe5CEcYFEld9Mfs18
ypZzPdeKK3GO9WIza2OoajbPvkNxFhnUPyRx3K008niBgGrQhAgzMnysv6vGsANyU3FZOWkv+jho
uPoOW/EHBuppNbVrLyM6boQedlEWjUdfEbxBtzQA+LFhqL4RW2Dc4RBsus55MbNeyJ0zXqgfc7V5
QYQEzAXI84O94ECTm1okmne3vxSy3KCKzh42BAmbW86asrQ/0rGRWTTU9FJamrW4h7Ksd+yGH1u+
VHO2lw++sKsHkqwLaR335sb+yu4gN7nYZFXL6V5B64QqXl2j5NwKrNCKp9YckSn+t4Z6MAe2a7r2
2KweL+8k8eytOclo/iTWdiu69gl4GXFY6vpM3OsWKXBkWBgTRVbnXK5URdBxy+BQ1z/z7sG7RFzC
FU3yfB8OenOOjsk3YplzP8HIsnIJjXxXTL+7KnyOdIxfGE88CHf9/Jwn8XvpNcymjQbUBDgo4kmX
4Gshbu8SkFYwToCd2G+cZ0YDQn2xD+UStjvcIh6ZuUk9JfzxnRBo95ulPekxSw531X4/Ppbw/yc1
7RUj6nuKsPc1OPpg5hBWkiO6KxVGSqSr4WOX6k+pqfV9z7Wm21TJw6udz5FR7P8gg0v5UF+TBff3
zB9GIu47Az6SKE1fXYngvx4ZixeQnsGS4oYut3QEJ7AZH8rfaAXmfzJqd64Q3qqr5OlKS8PlnfEr
s9zNnFfTDYxePjl49NOu7p/5/lT3Ycx6yVmFUxQPtR6wkxSYMZ6vAyigKK8tg4SJ9v+xlJftpEaF
4cA9sxCN3EEKO1XwKvyF6/y+AkS4r+xYTqCByfGuffESR2S+szQFSSwydyuz2YuxzEoQIPhFOmJc
4CqGDrGgMhciB0Cc1RyYwR42coqODiPLyncLerPlv4Sp5fmfxaNIUVH88s8+YrRYQ0MX38Aau3W1
Ts58Xfc/stUSX4XTdGyj2cZuSS4GNa1Kp4CBcA4FUN7S+wT1gWGN3p+qRNK6LmfkKJRGjNG+cMYA
bBaKeCaZVyqhligy/NXpxXWBNm8qLbDWru4B8sN05iQ+TxW842q/anUqpKFe8TpmrIqqhsN6O7pP
fo4lyWxnuzK+vViRdJY3EHs/W0N/5Cg56U7glfQAS2fiVuOc+waFYKIldP1qwVHAwqUbryAWhCym
rCvwlCmfc7r3IhACHgMR63iYRH0QDHLh0mgxKkqKYJ9ySU6tUMB3fM/gFUpZZErm4J3ZdoOjnicM
9SD2lv+f7D+0VTewMZucAcJikAhP2WB4L705crXNIA12magRaeewQc34P0Phe28oVOSoXcVpPuTx
gWvBo9l+gTiwzuHfuKn+HmJF4xFUn7i9nEtA/Dlwt6iHJoEX09vQt6RRmVcEab8FlBhC9RHpr/0f
TAqXLLHvnd7FgomIDFiVc5U2FQrhJ+nQLoZcW2kFqg7Pawin5OTSUkb49IF5DmTF/kiMU8mxC4ru
0a1abu+zFlvi5yyudNhqtZcLY/YAZfZrQswMap2kuTgLliFYhzzS/DgVdfp4e+iiwNr1sI3CNBdU
ED9PK9dUmZTdlwxScEC84djnnSKIjD4x6/CisM2qM++crxHRiYdFHZd1gkvcYAqXTwoM24YSVZrp
NcSdxxcv4ID7K9lNuG19eztoKC1Aeo/A3tpxwCRBi7c7zBbjlM8TPvOHLLAJmcYK+mv4TQyRSXQ/
PwQfKLGOKIRMFR0Z5/9SDoD8dLPHjs250j7a6YGrbZYjZee5J1idE+7fLfZ4AOuUgj9wLn8IO09B
8VAq2mPFOAt/JMJY1ehEFcXK8dnvXQVQcSeLid23hGZsANMnWBdR7Se5sZJclFwfCAIg4MN/k2J6
AcT5vMEhKMMiA2WPKFKmjacXiPfrGsHQrolN4m2+m3ima7AvnqfvZhUFWVRv8A9DQHR/q/AfHrci
TpyToAE/hut6N+/BEP8rIWTfKNYEmOCtVxU66xH1o4JZW59Rj7a/jHdiSXa6MuohUg/qrlgpykdc
ZOD7cDL2SL5kT/LH0cG/ECrvgdP5vxY0O0MrH2EP/PjBB0j+NXOTtEc7ZfHpMWhU67iaq040qA/x
PzFpGdwOeVJhOnkupN5CsBgoGKUqUHouSbb5CwWc8o12M6kKA2or4tKH6v4txFPOjIbg7+7/8KkM
vxxfgh6YUkmBGrEG3dTfDC5gV0Of2jQhHgVjaX6vJ5aW/jc02WsbX0yAfUhnK9rg91K2tVTsuRVb
MQ8H5lxoTCLE/meokMVadFihqtqkPw53cCxd2gYIpSYgjZiMxF3KTh3/TvFFojBq9kFHqrRS1Xc1
F0fxImlXgSBAnBkllOp+566AvHklsvdPyhFFaH/d3hdnnScDGyTFBMwyzzLTto/MngdV0UF0hH7q
4HwauGY4oYtAa0mrXN9G5Kq6UW0Hu1xXaEdBqksWc30m7gBVPj9c3+8XBRufu3br1z0tZAIr8rCE
XmGOupuZsbwP1TyTSmQx7lTap1dpcSBHQXqpLD+4K5fEoi2DvnMdtJjmxYOzEKCQKRXyaCci898a
yIdCa+iMgfyqc9pqqfqKhedkafHGbvSp8/o2nomAtTGu8UE78/019mVw4JdCn6o4c6+tagLb7LlO
pQvjtH6ssX7MqB3xlZvKEsrB+u3CJBivz7esEASkElPx1jq1Qw1vgBNqNfVL8gIhm8KRoa+DrLet
xK/bOyIVEyfAqDQYkuso05BucuWKeWbH2aeSTEeoG8Nk35StndJUmfeQwDCxy2/fZwu0FMfiis2F
8JS0hP70eLET+tEu1SvA3FXf4rD+ABa4fAR3XzRBTKkRkxUyn8XYYDX9KNTk/PLxVBbLwHBlA4ht
UID3hjCLSdyyKtB/LbsN97vXoIju0k6ideuBgXXu/oxIFMKGBL1tze5sSY40rNjLqOX2S308fjQ+
pcYoYpugPBZ8U3kY7bAY1pzE/ChJKwdZI4vify9KTP17NEsS0TNfvE3u8Vw52suXFrL0WisVHTdH
DLw3QbfUh4PltHdKGdgyW0pMB4N6zYgfoEd84pvn+Da7JoSF7YaBFi4haHfRCodN+JNGH+OYx9Da
jJMo1o4RKdNc81F3bHNwcMF0zkfl5J+q+vqhtahFEmBYNv59HCkrsYOznxP135jRpgePUAoMrdAJ
TTUbixB6Gi5pmNJGd8khhOF7ooXLbe70waZV1xIPe0m/gfWUH8JN24k/kINHNiU56XDPgxXLVRPS
1wrivNQoL+t7lGXeQFzV9en8VBQnDLkuFsfRZXyse0mwQLU8srZxgrp58Z2G7Lld3pveKDqo35Cx
XHqugsbLyQSrKRq3JRPFt4eyTfD7rDksae0BYR0xEHPQ9YD4ntif3nNUv8MrV9LV3CKmyYeHftCW
cMGKKcOY1aHLn8WSKPE18cI6FNE3LqW3Ctok1sKhmfHChwiKdotItBFd+foVi9qfG/oAGvqI/PsX
TQmvStJqQ8qm4fSOGadFvC3gy+2arYzLvsFl2kRZGmwhbUQ7ZGndxm4XcQjrlf8dvjJvDB2uC6M1
couk3Hp986f3k+Kc7NFEB0GNbjCPudd8kJ5R9E/VNd5mfhMSKJb/fiizTZy0KFSrG/+SiLrCjIGx
aY6FK8D5dutfrkiqo/dGnKZY3tRNUNlSPld2ApCGoMbFNUZyAB2xAi6/yLtymjrQbEUIK8nG4G6+
3Gnw43z9qaI9vLe9K4OrDd6a2hkIrOrKaBe2BD5JwGgqfu+sGcnxuS2MxjREyla9//J/1JHOLzoP
sB1M+JoIE5GL/VZMfqmwH4hBeJqJQdX8j+AqJqJSDdCIc5FveDCfEeGTN83A9ne/ls00CwOs5hmx
UPfLtW2lTGrKe43YAlXMIaZaAyKbLUI/ml16TBF1OwJcpKhFdajeEl5Z3iEqb0xS3gLJpRcvjPYe
45hm1oQLY0nieTVrk9Aim7vzhkW02D/5BKvgL8RxTkDuDHOtX2t4LcHNdMZSW9FPyD7p6X6Y5JlL
u2wwtdkKOhYqrsWksza2rr2tP7hua8/ogihZI0k+dT0kxXxnbLo/663ebkyk/1d/K0RnMy9ZK5Vh
3jHAZqBaikkRCXLv+S8nxDPb8tUqtR61JmUOzcY6EOZCzj/dueDwhHzZP1tC28wsdg+2BDPvO0J6
wFeMzsIPdI/MCMczBmzoQo6w8y/iv241FN5cMCW5huQHbXOSIB/UwqUQTCgybYolEYV9uiOZNxRe
wJrYbk4PCFtB0T/ux6gnSe9zwvseJFSD+rtK3FURl4wCvABhX1VtZ+wcCNDyWjaBQmatu8oDSlHY
qSUzirritbNPAz8JkqLoUF0OCwfBo66mZV5hzUUYmAaI8beMabmnId6KNz/MA5TlDFY/gEhG6ArT
1HE5ciaTg0EwxMacmflktSq2Ue52NAzDsRhTQxBFH4Ec/uQhheAVoT9sNQ5cDTsbP9mMFBTW9/VO
MLFGzaZgftsBxZKPBHMUU1Jgg87CN+pw72s5knr5XLUkgG1PbrJLdNBg/0S2Cv87ZE7AFyyJzX+C
E7GMfj+q6+grYL+EirHb9St7L/JGSxZ11NDWeuzDAPfUxI9Sz/IIQGzZGpNqBHZli+2kZHZ0WTck
o1mkECQxxmKpUH/QfGPByU3/SUoGT9L8mxDsvAg+u2qrW5JR13OrZWo/vl9ZssqseIRxIz//h9At
gQjM3qHkKYhA1yGjLiCikDiLhKeZn6NZTwqD3w2xjZs/QEZUiuaZ8Ex2wq22mfpVNE4UatUdNlUm
ldDmF78QaM209P8rT8LzcraTokUXLEQ19Amsfthwkr6TJS5El2SJVrbPTrY1oaJ5W/SgsOtQzzp+
rkzNbHY+lEXCnSDOps+3MZnk8FvuFGK0LLCi81tt4241FS0Fun391aDr42PNXQ6VTXuxL1/qvsLQ
Ra3qcmhoT2W+ZO32rJkHARvRNis9xYTjh9SNJ8e8fOUSbVae1HWks6UrVcUl2E0GRlxItju4FTFJ
rjOpw1Lo8vpvNV/dLdk2J9GX2Pho7YU3ZeV9E+NmyZ/m3UnVFORz0rflAfStDiAHovEcEqtW8WGM
qOY7WK4JF+30B0PVXxxzMTM+S9+On22uxve1A+BqmMpkdBsJYBTcmQKENuDRZr6Y7ihmQty2qpXn
Dk5HsIQvIozll9fIfuMF0t9mVpd3SpOY302cX/aS7I8ynZ1TbaIt+7NgBd61A3vuAHlWl+MfIIkq
rHMhM5/ETwW70jnEX0w/GzB3Kl02KHvVKbvPs6KIIcWCf8FBtBTY0nnX26PF/xmpwv2fqruGvbPr
4/hbXSv6s+zLE9remUYrPBqvtSXtCFEHmUBmWCr4ZTe3JJzY7FwgcMi4TJO8vJWl4QWuYYpfUnK4
J1uS+dSHgTAzIsT3fmBpFfCZB1+0OZ+PUlLsCoEvXWURuwnvOTWPxfdJgT4r4mgvm9I6gyocPNiU
W7NdEzCB8rZRfLCK7PYbcIHxrTzIGwXL9E1k0SHOGvoxHErjyCIJG6VrupsFD6fxc08yUHmlYi7d
2BZIBkZOGNZIXqguTaFa+ezNN+qeZPBzJz4Gl+2rK/H7xxZpYZolMfEWQzaMGAkOmyiAzdif71kW
+4kkZPOo6wR+BhMiev8nHKXz01GrsxiLeQ41VxpzDKlrfELXODTaJ5j1Yyn/dR0RYTNmaKw09u/Y
r0dc8F3tT3NLSeJXA+BpX8cgkhBNn61RzHfQrWjjv1K8rE0/hBrgxosMT+S2rQKH0BBYiOcp1gfQ
IYudhWPQ4Bl2VUSKXxufAKf8sVm9n33JaAcBR7CYXrir2BO2N8FUi4FKMKRS8/ELHbkzHbFbEXi7
ibL5eYrmIwDN86kWyV+e77l6ACAJ68B8txd4JK0wG1j/xjFA7ucwwLmLQQLyAE30ukVIXrtmonNE
Mc/K5PtJXF9jIuy9VcT1jYAsi5/TQ776yMO7HutNxwjriiDvRjsivwRkBBcQ6yyHmCzZD6i17XVY
qrtDbcWU8cm/hQuykF3PhebSzBCKbuKF9ZIirH7gXSnvx8GUONhJsoo56Ro8QTkNYaw/PuuwobKT
x6/JCxhRyn63pyxWD6vKPMP/+WGAjBcgyDsMEmKNP/yu1jqDviDAk6q7mCOJNYA7ahJOCSxXFEfp
3thM3hrvsBZzOuNxpUODgjNLzfvN6InMuYOI1AV7JN/NMPx8yT53sTwSzAFkinURUeENRbaDirL+
LBEmboSTgNurLmnbQNoEBdRgLMV70y6wAVr0CKg0611+WSbGhk2k2s74eqsNAXG9D7m1L3soMqpf
QBnSR29bxaCIvORyNGzE18sWkHIU32nTETzmMAQoYlAmnSdlfmdyhFTE9UcsLX2kxpMO8+XbPtXe
hIGd6TmJqEJ8p51ugaDSu79WvGpiBPJLKebTCc5VXpBLMfQL0sUpiy5C+mjEh97jcgGKiSg8AXJe
3Fug75RBsw4k37TqqDfwT31Kg/cqrJ48sojzQJ6AdgW1Es/cd6PJHMp+JgD+mNyuxQ4heylDgzpx
81Pqh7KPRDf4CKmr09VkHM7S7x9BGCckBP0/KtKCxm96r2DnGs6HphqeD473vB50KeJG89x3WUJJ
4RUftZpbSMQuRNP+OHOfBZ6LkiLtjYPbd6/RPAz2jKbW+9PBpLO6qnWSrBSp3ABew1/kdot/v/uW
GHyyLEBaxokbuE7Fwp7baxDVyfA5qNHD2zbEH7HLJREjYNa6CzIY5DuGdbVEauZhgsXxatizjvS/
gFQq+3JnTI247c/CXexeULzRFW7CuzJg1x1cQ6ZulXltC+eme8lfoeNFozSXDTHkudtEMJ2zkXqV
CGrSz/pzaWTzvHKOomgU/PN0crvmalBWnVfvQY49Ycop8VLvJcrTqJba6da+hDoM5ClVVe6lM02W
kECApeoA0w9r2IGf3vi/73bG4QEA09NnaUTPKq3FprWjbZSWVuo0JdOGoN/hkMqutbf2DzCfIRyi
q8WCnvNZ7K+agqsTXzSQaE/MlWBzoduwdJtp3p6drHGD6i2IKntTwXpvm59EbkcW7z8Obxh0ILEN
g3lrcsPQwhKgEO8pP76Jm87lgCxR69j0w1rg0VsweOW88XdmUhxkKYWQJHEd9x3v3YenEnottV6o
q+ybKdAnid91QW+VvJh/8JwdQxjNe9d48Cwb0G7fpnky8PUOpzxG29aj3KZ+0+sxfkrLvCrw25FO
geb20uJzCBzw9Dv6vDOXAZclTK844ISsIfD+IVAtZ44OGJZQHhn57jqzFdxu79MM0dIOpDk84kR1
8BDb9agGbcjXW7JLXXWC7eq8qS3UmLVHMpDHxYbEDg4lm+REVfkAbMbkrw2zLdBo3t0vlmx4vGtj
jDtOgENJJdGkbMF2oVZGwe1/0M7y4kj7LtB0/Fv8kUhn8usuJIuamTeohJcD/6CBVKOS/g5/V5FH
exeaspmr57WT+CZOj3S33AK8YKqG7kW0snO9vAZ5jdlJGC3oqtJatTdE43Og20NtlZsnmiDVGfMk
K1iYty9rdA2l+E5d8J7M/b0W7BQFajX1Wphx4kzs0n87G2JrBfLPTgePGcE6WXVvbUF7f6hb9MzT
Y6dL/uygdPnUl028VdAEgDYq8jDrJflxGv7HgwX1BQU/s3uYicgr148kUqcF3E4kUYLYBsUVGRZA
2LEKKEElbrPtU21o2IIrfzC6Ps2hKHZlpjMGm3ClcRhwCixMxM5j1749jiLxrssy9kx+c54vBtEG
jj63sz6xjHQWTpDFhH6r7fEAph6hbce4tMgSE//QGJgLPnjCQH1nncnZgVHKdIlSx57aP+L3z3Hf
ZheQ9KR/o1PmhF8F4vqD0M6w+hf58gLN6Zhe76eYPsWaDHOrwAFz0YS6sVPnm4upqsXP1DLj3GQm
+YroF8jg11e8RtgSqwgwoAruThLzNCYk3xaC9kgBzw7/RRIXxGI28Z5QHUFPiU8p4v/5iI/0CNbq
TyVblczN9yzG0NHK6jwz65te/JFIGo9dvbqEZFDS2aoLKGKH4UCJQcgsAiF1Ixntuvo+tHw+7BIt
5z2fglt5h3ZscpYKRINmaNQjiGCyXrZzFrh1wAmCPdYeMSyE5Zu2Z2XH9VhbiVxOFJulqVcx9jB1
PMBXZ+wKnbqx8ac3ai2bCPLbez4MQXoJvBBUdSG5F26jTfg5/GcGYwsYwDHV1pD9T9x+3Nbzi++f
yMZDPyaysTiPrAeJ0ujdJY7Pvt0wCv7Y9O3K/e2764GMJqSi45epS0GVLMXfUMS5JkCVGtkKJXZQ
AbDluX3wfpgES7xHgpIAk2Yt1SUAdlI/zEjnqdsXF8PSJXt19fyYn6pSJH8WEctxAyQVWUiOv7Z7
6IkYTRhT8qnKJ5YwOfWoRcWBfe/YCbmLWRFdDsgyaGIqOQgrUuwG3Y0p4PBhYLjS3YWYramdhlev
/rJ65QuYnFr1wVsa295ARyaxUdeO9Tmw9oCHIpUeanxZfoZP9sd1FBhJ82rAiETG/aDA6o1iGzTs
kcn12l8Xk0A8BuCa8qJgm8o6rNj8nt4hWf60+NolOH7XVnMLrDZ3x8f14LPXIoq7AuHrljbXqEdO
YFao93HjeTwteeb4nktr/HSOqKMDtTDfyHS55Sd6Y5i/dqrKTF+pw/Hl3TFZJpQkYSg3I8uVGa9R
n4dO+uKNIxfJj3Ts3wPTc2BLT+lORMtVBjYV9V5ValjwphP3T/ROnyUjBH0BzBQ64RBFE+lQrUox
/7PpYaGKqIgLZEoqmdpLq2akYMEuQm+j94opvfyObI7wOqxEzD5pXRktMoQrTCToLx8ff/x6Z/qg
RS0w5K4VDQedqB8X5w9YLpxlCP0/UY/rUJy7DeJWev9W83W5yE7+OVbtYyluKsPpeYFmH8Fr0C/e
PN/Xtgg9wGHot1LnI7lYge/JYL1hVXKs/sh+4xl6byNixHfSs2P+iNMJwI7hIFOAoF7OPWZKejXN
HL/xskQBEEG4dPJUuqqbSIP8r7OcbCJZy59zJvB5FZJezc9soMbsYkuP0E//ofdK1fO7iZy6yJ/N
2WUa9M5Ks5Rz8JarubstutW5mU2/dRoIlNb90Cs9aWbi8kcA3DiYfcF8XfdYotJaTaLWE9G2d8Kv
ZXjGUS56DOts1pdPHQq8w88lqdno4BDVSw+vrFAtRvayKInYFqSoGuTHXQkyUcHoxDfmn74qC6gn
Nl8ch9LMQ3WYdoupTbfp/h1f/XotUy4xLksC2bisDHGiEoOHNoHw2No4xjVWDEDHJEGNtPVc4sAs
E7VIAWGfVaudVEBgwCFkwdQQ2zk8juryAJI05kxX/2HirMaNH5W0dyD2mXN3RcY6PqYKxWhJk+5w
7y6i10Pu/KUB1j9ONmoX0pZmlhM+Bj5XmE5PmbyzjlF1In5z7UuOo/uRj/AkVmFP5BS7WSUJXWbB
O1XRWHZkQWEFG4htOciGkNaJPYaKy6NOdveH+8XhwxZnYJPyPi5KV/TsHK3d+hBYWVJ350DleLUW
II3/RoHgKXlmvpFzPtMyJC1l+RJ6Qbp88eEIbVpk7H1aUHA8mIcJ8RjTOvDcRvalI0FQ1HeaO0vh
+B9SGT62YvbZR8xBhDG+uK//Ya+bBxsoS0wEWm19089JBpeX0ctWzXOcFsN5CJoP2XP8rjDFcrkW
HPqMVKTZLCSI4hxb4VZLqampOtt0eaJphvM50d/kqGShLvhzetelZS2xmAbqI7WlDiRHA+Fu5iuo
Zdpojt6KR0jSTf6lDip+sT8z0f1ap+OZKP6g5g8172IvH8IP7pQpy6AOHgcrfQ5CEzo7aFUxgAMn
7A1Mo7dT44kLEGrXlxvN1V3trY4du9zbbiwQx9KsAKHDno4GymMoLW4t13YFN+NasbmbTz1SVyM9
0iRB+ZseGHlmfBIwuZKbUp6R/z+L4+6XqM3KGs70cOXS2qDagN8DHRWT9+xk02Y5PBz4Pj77mJEZ
sXKjlwPsYusEQF15x+xWaYxV+pfbA6+xlseS3zu2yWFiEd9GjJGPJuuYvFjEmzEdLS9BqJmMNE+G
PDoZEl9VkPW+n3rniGLXyiDL2Dj1AuTTLUMrEYqXKDDHSB2sq7SPzKbrvj4IqOCUHP8LXnR7DVdW
zljAq7G+yPs4C4ThYaimmp4vzVpJCvYTpKx9yGaUiTZzsvlIAdb4Q1GgCvbVRV667rGHVi9QtVe4
xClqZDD8U5skGr0MZM+2JzWdJZ9cypd3EI5+t6V3EsNE7/GUNVrgkDhhtUzJnGFUBtgG6/PBR2l7
BLvkbiNgqmYx8OBLL1clZUePNcGI7BGAbzg3/vwNkG3gmGgxR2r9Rg9HNMO2Odho78QNjqCzx2eJ
2aldBi5lTK/D79razvqhkaOT3mOtP9Uuv3k2TONHNRXLbDgx/VzMGwKJmp00GqwOGg4MBzmVs2fB
OhVBNf56CVUk5w+6mI/xz/Uex10m4LPsCD1gOOrmYSlCYfYUu0yMyls/S2T0+yVR7up3oNfvNxyZ
eT4jbDjNPKx8w2PqA6wPFMwGwgoPIkcFU6NZFXl+/B74jv58XTeBhT/P+4jWigg4y00XMR/bYkBm
BV3d217Tn6WjQAWsaU03azKbH/4kzkW59QyYpv+RDlG2gkl5euwL6GWC07pV6kkIi4z0fKenhwPn
5c+pgQY0Ts5sdq5MH6gAz/FWmFOY3eKJYqW9LlqYBQAfcJ7mCue1b5bkJjCSvLGs0x5/fOoOIMos
KQRVmtQWQCU28KPBAuyh2vZ+jZXpF11/BAKpaWNGOgLRjSf09yRuBmv/Nl0103L8nXSiId4HTFXE
KL59F9UhmIKHmDz965cy+1Hhkwbq/2IGZa9C5mSv6kEXKNKvbcitleVz8I06PepkxUeKChRpwKwV
GZQ401EfwiwTW/ANdsTtHH1MwGGks66PP6/f/CgvLOgxN6X+4AVc6nyXbEIzR2uq1Pic6+IfGPs5
DKObRoCk8iW9LKYbfQzq803WCaeSssUv7cmJ+l3Wz0fLH8pkkC+IFG7fpYo7F5k4V/nnZc0sPPmi
qKIWLNgIlzxIxj2eYl96TOuLJtyvIj4qba1DaYR6KtMdkcOFtlmAi0b1F7cHeuTy7qMp0FXBGj27
cixNB1UrxY5JnsxRAoqRsJuRlZ9Dmb5mmmZfYTarrQACgdOPgrgRyRYx0zZzvPcP999GDYEq5aDB
J6edEfYxpJibzqCySmuM3N5rM4JHFNtYxgUZ1qu5zeWh3kqXg3szqZP7wKCwHl1c2zWtG2NHtPSP
qp+lcjK6ncgTmwoAJCY+sQEk/GKjCMxCLflFBpu9lRwVT1GDq4iK+OZZwLJtN/dz5wk1jWjdJFQG
Nirddlp+YSvjRtv0Qt7ZTsl27Y1bl+QbnWuAiH6fatuU8AzUAEaqYWtg2c0fdAChDuXHWBDVoLIx
4h5u7B8q0F3XY+sbohKxJnsocflNV6ye+IhC8HGL2XuhLgV3VTL5iGdaqc+Jqjm1X8x/qhfsmEMv
Y6vdQsSmUSHYYRW16YOi6hftIu8UuQOeMz9Sky6eOmzhKpZdEnfZ3JvOKMDYZV8SmisLkC+d0q1I
L0RBmR+wHF8FRUXrOerEHx07rLqF/iAKqadHHP55Q4jwklUp19d2/SC5+LCk1jldN1dsQ9iyk8zA
9kt2FdY1dZgdGfVJbCHfVVOW7j79oTJ1T/NRUGXUM68Ug5pSaeF7K0yTm7Nxy+q9lErUHPmsrV2Y
aLCj3uq+0ZiiKDWEHZ5+OwMd2Ack08MHIoVPmaoMWPdJWUnEMHqHs2/NePC3LTZZue67JL4i3J3s
DVbp+FBj4tE/uDGUpvzeVFT/T2PGRGZNcXsIZUru1+ckWkcAohvlX4F1WHQd8le8pBSapa6u+k0K
17C7YdoBBMuBRCrT1Sc8NQgh7jABHe+6YKkeYJLEX5xl4xXD5odzEekIqjhUk19nh+BVnPn9DuTM
Q1uhtd7q3GpPyXZsROJ6rRJ2IhVGExzCvlzrv8Wu6s+WXcXYCDdywsSh+cU/DHmURjUB1WciNXiW
LKTmi7RLS8NfJI5noSmW+fsvMDhbvgWB6oQPK8oncY8smUZ4OUiWOhFn4b+psjPYiKgcE509ui7Y
gM0ZmIyyHMeV3LZJJpCqW6eb9jcAM1k/3nIlPulhi5uug6Lzd+WNYV7Kf6oef9EATQ65dXWXbqoi
8rDO8QSblIDvX76PWnZoXSN3GK0PBXHsU5NoTcVPAGIZHMsRMyLyvM5zo2+IbPP1sfl3+Qo7Ifl1
q2Ks0x864VHbWoOmw+8sJ0tqfPtYTfTOfBTBgx1ZVGq/ZTLnvRbDP/SUHv6cPnqBFBgyO6n1GJZL
XBhXsqgJRoBiTs6FvUHrq4HtqGkUyTjrx7biMEyHImYx7d4JyqKlDcIEgl6TozXZtA/NQOuqn9fd
TIPx97L5311nw4Rd56U3QvTpZ3yLa1EGJUKF30+mR3oZcB73Ar0gR46hN0b8+fkyl9ETfKaoV24n
aP6iMAie+DyQoYD5l3CqUpOG7zU/OkumNotH0ft0mrj0xgsTDw7YIi3nu6LdDWC6b/rdxZYXKysK
/s31aukQckUKvuPmRB0F+MAUtmb0ytdqQgHAHujqzO/TYOHyKTu8Qtc/GR9Jp1Bybk3EoxdnKvWE
EHMppEJEGW5cq2C/OvaQ55G8WmFnHXghE0HQvQUJee2IxrgmRMV2Z8mdypp0JLCQcGaH+xvXYzLO
51q0BB1iAltY/Z6o2wyY2cmoSEuouoTflQhKBStjgcsPGy+0kjGny4pL/0vLjsUNswobATd5Wa4o
BaVOU3zPcgCtwDPScdx1T3plD72ifzp1Qgzuhsd44BGvg1JeLFCT2upyLHKjthlgdKfEXH6ub5du
kEObEBskgurDI2xtX7epPfRRwwuPtGZFhU31IOAWyErPDMW5vHcEBl/cnLJge2BzUhyOj3PwsOxp
hFqmpxGPQxCMaOLITTimFU/+c4Tg+bxHxB+vPPnr8kNUiszR3Tv1KNxwWwmfKPM3MkMekQDkddip
TJ6vD3K8mQuMP94/8MsSOXdt1Shr9aNGaRhknWKaT3eqvrYZU8QiIBMW+mx3QvCBT1/1f0AAPLfO
ht1TegtmJGg4bgygLGZ/x/PNQVSgrV7/2k31oAIaaqU9nmHRPCv7gDxE+CXqhr4Iu85AZdTf6XZE
+sEjIHrTskSTsPqu4jfdcxST+Iad7pAT3PMVP042m0niXFdmDW2Xp9pGTGby/IOQcT//Nkh4dEfS
xiNhriOZc+to+vfkMuYaIozE0KyqxkJLvTydwFTwLVk38mbaW/cig+ElFwGLZMz7rONL3szucNNz
n05JXy2CfctBxWlj3hfyeBOvegIklJ20WxPdClMHNGwq79ffzqm777iu0b8SMTt8KABW7bYm6HDo
88zfISVBq2NCANXFNDl1/9NR6ZSPkYc9xd23sL92+a/O3llmnDbHV/EmidF7nkCnnvCqnw9rgyWo
IC2ThtgdOGIgdAL7jKBzKfrD2wfNhbYIIuDlUrODsNZVG/cyIcHoaDzVv91k8NBtSaIKaxfou+kX
w5oh55p2+L++EfEt0hZY7I8r8nD/AKLtWAJdMR+PSj7WtgJm7Lno9J6gWa5b8LFNPcJeLe8QiA7t
JHORo5H4vE9Yf3Uxi2rBY/cpMA0CO69vPpyUDJ/TMX5b7oFSYYMpdn5MzAxlI0SCiA87SO565Y7q
N1rtqJlGnVUlgAJcXHxcaXDAClgx/h9l37k+WXNDLfA4f6KSwicukqKnsJiLbeKwKZ0Xg52t6vIN
jSUYLc8l3vA/+xNDIzsPoNH6J+BBb/SPitG482+3udAfTjTVXj+WmSlk/ubuER1SZjp0yivQzOo6
DC97UGbRl9Ha/OhDODAOXLluDkY0YIC5crgmvZNjO2Fc4bKryWR17w3mRSzclf94CIBhmSJZ+dza
mJuudIiLzpYFt4jszinaLRmLKAvrM7yJedpMX1KPoFffOdoLZcYWWi1dbx0V3ecgPg0k6IRnDQsu
8iOvXv06Ms6zL/F9T2PbYQmDKdM90bwuf4ICvkNdRovZf8YiT9f8bwS03eUYVMswL4XCYic7wXHr
LRNeqcZmZviLtQD6vyvp03LfhC58upV9bnnpuGu9q6eX+wvYvx9JBfL/q9x11fwi8LQRxvra0MAz
ulG12BX5NaAFWgseok3VjlWSLRGSIiXKKzx5s3Temu2sS1mC8T7p/KmDw3qK7FN6tpeTykfZdNH/
ht0vmqwnT7cV3EeZ3yh61FdkmcvqsX8vg5qORpdfBDcJoIqMcJMDxHPJvJ7gH1ZIs2w6qnlcVV9s
t3Il0yONOL89/yGixsMXq0sCNKp+gI2NGoRZs03MMSW4TXaTIRycC99qBKfi3DMQ1eR1Ls4ZTr8M
mJLfmLFU+91oDjsn0LBJIWl/HABCGdwWImzXeoa7wSaonjhnWqAHpDwAdRirA8uAkZ4Hh79KuRCg
eNElz5mcVqGmZLZG0+ekp+uQijZ/Bj8ODJA2B8MqhydJNIv2tXleImFkDGNhvAKgRATn5BWtn7gR
/rRx+Ia/yWAaMNT0oyYtX2LSeRe+g8N063ctNM1QHwtm9EWmhq6dX54gVq9wVVizew4SHjd8EizJ
kUkTrinxa7gPX2usAZe1Q72gG7F0DQBA0UBK7YlDZ6VDoi3vn/GXGQ14sLX9qRCVoOOrGnjgrK2F
yAFUCmAH7H98jU3avHib+QD/Dx7KpFrLrPei4ymisGMMmqfEhkEytfG6Dl+IYeLK9rRMtRhs0eZr
9auUNAP89fO6/RlhSGOzuyYRLCJgbhWjFvof19+J9XQbAIBvs/sFhgbpLq07jBjrVTjmHDr+p3WQ
WNGkM7u2Q1CmP4FlMullxUKe641DYec1hzm6jpRr03ESkV3rj+5PgmP6uGIeGFPCao5bbLJXFkgk
fik7MaiDWl3YCRWDWLqePac6qzTLNaF5KX2RAK/SwbpW4oLwseltrYuWmbpNH7EbiNTW7UFDxinZ
9gun1uBJiqyjnCM9ckPsVYJdbJYRb+QoKeQM4TzkUMWE13ukq7i1JgY7AUtqL2+DGFVq6NBNmwDH
4z7WfK+pfPOBJ16NBl/fG0b9TgEY7vO2pU5W8bGkstKBUwzKDPsa1j7Q8PX2pkwhDiauDAu0tkhF
lnErtOeDdvy099uZ7H72C2n2Kq2noe+8NS32ACU0fcA/E92Jr9IEDXXNhpmDtrhJpLRjqUx6O8CY
ZufUZBUZmiBpUqJufe96FHMRUZJtc8MVama5lBqMtOrlUOeutaU6w86I6hbERL/epVIQ2Eh1UZyb
wgwRLMXGyXZLOEbqnKEGYhj6aenx8l58ECP27kC98N9J+HOnaW5ppN+8b8cwkxPZmpZZZD9Jt5Xs
ftWzVXKlm8Po22ATUafloiA5+RE0nNTWco74BhfUOBgv78NRyj+nswIM6Rp4460yR+zbPcMGJDM+
RfUXENGjWRo2mQF6RYhOrtVWVGswRAK875U/2N7R4lnVUfX0xEaqvyVqHYEBwgEYCbquNJ7fME7a
708BXB0hcxWN99uWsTO7oCamRqjQk+6FtythC+4AEuxQhpHcOy5Km7hOVnpcQbTTzpMHjkPt+Cz2
13jtgjCkXsVi1ejsVjuD2qs2qh+uJgAzl87CECMaDt76x37MUV5D3OyDAlNwy8cPwhVEidhBUSNa
3xWmOXZmWbEYCV4B/n8M9R8ZsO2CgDVfJPm/B67rLrjKa+GMZ2TuiXCC7p0p2sBPDqM8RLUlYHj/
5XmNMBbGENk/9TeVBOmQyy7IsVOjh8SwEXs0BaoB/Hwy+VFcXx67oILZwA+0oUX8jseJHjM7utIf
Fcb5UH35+WiuQjeag/bNKB2kz/uKJ4Wyc/pVgH1oq3vLgHMA7/bIB2PzQ4X51OCHWsHpKNgkq0ue
QGnLbrmUsgInQ/c0H2wCfWJyWPwwmVG0mwHlNQpzeirpF7nosqLVqFCTB9zqapsjrjXMKp4G1Lxr
g9PQyMYur9RO9n0kquWBI85pX7XvH1+vMkOe+MQeS1Qr4eT2jeWHCx13u6TNphA0wtFcnDp9Qgcd
foRQRgdeYBoKJvcLD0eJz3OojhLdL9EmvW9p2Hv4ehYfDeRQgNSyxYCMQnxUfcitU0HzfsB9HKoI
f2AsDpPgKzoT/kwdzE6qEguw+Q4x8zgp4rSolHC8e0fNzmbZ39MhTMr7L86D9oY855OV/A3Ivsyp
btekOuC7+ja+oSDv/rRwlV5IdIl3pRdj0Qvrvo9bG+o8N4/y2Uasx1TrprI/XgKhDIyY89HP0flg
1NoHQgJBnfCTVtys3Dg4vH35juMyCfiWF0rzB0SmYFMoFDLHrXtt+tQg0wsHX83abpXVNzjqYBc8
ULImolUr4OiWK3E7T9P8AVSs9gTnDUX0CXGkbCqCZ2uKbTAtJaGeok3vs5Kvc/IB/TrcgRVZG67v
Yyn1wcKphe9o4coGw/X9zmimKCBTya7k4Zrl+Oe9fc7Ltk07REUcgQL0o9KvR7Wsk0GswOveT7kr
Q9++4l6TD7rvMpVaaRfkm8B0nQdOksMgRObeWTBFF/mprJRSqBMNRXiqWljiJyzwVRyLQGBjb1iK
qX7OKqDuuZTSv30AZjUBOGor/hikMV5jCaBRvCjDUC3DyFfOB/pdCGPtFh244hGVvrnz2U6ZScVl
WLytxmiTjMjR7B4j4IRNTR2nalvUS3RuVy7H0uybPI2ubGitRl7DkeJr+NmCz4aFRnZ7BbVO+RfT
39tdkDBe81yXE8Tz4Bux54b/oFDhVRYP2jDi7fnbvlyM2BLf3E+SEWTaM2Q+EpSUKkvKyNzCYsVV
+EW2X/Wj7sARGejT1tWcmBOIt+C/XpCoej9+ZPqLWgmI+HRG7jgcpA2YZfa62p9r62XH9KeGSPu3
KtcaAsGv7KguliPPEj1jsdLbxB3IL8eBlIRH9l94CJjCFx2wJzHFldMq50S9i6ozYS7cfMUBT2fE
/mjqbYLtMi0VRMSuq5K2s8zo6HyiwZ5/zpl+zmeXzTTzOtV7jzzB/RSuY86ZcL9o3GTaXpURkX7x
pp7kUvx8XQIXRRuytdOi6VIYi9T8DTx3/zyGPfzyDgfKmSCIkhKwDP/+szHDO+Es3TOSSWw8w74F
QkoJRgf/ruBHsZRLm7nlCeCYeXsWmTdYIVwy0GnTw/TpdseHrtCrR4odW30WJTqzcU2cOchRdRHL
kwxphFrSkek68s7m5cqmWF7JwwF8v3dZYjBhyGlAbU6HNPxwFEzI725r/8FIl2rQWd2jfqFzy6mK
Jyr1lzQFN+qSJRD1xKSZ0waWHUgteIgyko3siYTgT1XDx0CVdc2V6KdDaEVmNLuI273g7L2QVeW4
65VxbODUu60mNCgjQY/LUJm9AA8w9/oSLB7dsp+/zz/zsp3f1Ehg+NMV6yDWGJYfXaphoO67yqSa
y8c70EaBzaumZSrD+uAgEW4auaSVvL2apT7IB/bHDdmn7lWKg0nFOQRM/UBj5tZJCo5azTCLyB5t
HlQVydUaqJrC3dGdSCTAfN6l/uNs6lqfY9rvYK4MxjHTzLOKj0QGPvbOwDYGCOimTZ2uOL0F50Pb
kmpepTi5t6JQOIb8Lp2KiLx1aJenp2aGvJmxlboxaDqxw5znedZ+qxn6xocxzzjsJmdGzFW0LXqn
/QpfBQk8ihTmRCjX2cXBHkz2kIZ65RAULff6ldPOxejNB/nV3g5tfIFa7p5vN8oqdHBUyVdn3A/z
QJMKf9VoYlUHlcWsM9bXgSn6Vhch4bC9Xcd6OgFVDO8ObNsLh5gcGbuxwcIwfPFYbp/c4EmpQHr0
1DqPR2SndvTngIQvd4IcmdO2RvXSTG3waRBJJ23sJDHQ+cL3n1WAVee2yRYRy8VjbQ/pASZvFd/1
WuBXmahiFXvtIB8aSOvORHqRfHVJ50uoIfplk88PYLhrW5gGgSirYYLI+dzcCWlFzwgWeLqJfUSj
SUP/nBNzgEEd8PpDiD+Dp4MPZN2SadkFKPod+JOz9rgBcVQEzBFTKWPlcJeUQvlTg/oFM0j4VmL2
9Bbqn2Kap2fItmZoP8fkHs94fW3weGmoJyJuTcpGmifSQNyUCsG4AKEGtqx+95nV2Hl7ZnuTJgAk
/ponouC4pdOEZgco43Luw/WieYDdA+J5du64XXaiuE9paBtoaBt844Ck3nbPrzMJb99v2OzocWR/
bV5OB4T44h+b/Yjl4dJGbC+fSD5JkgHxg8r/fAPMnsrWipVj+/XHa1Yc3ihz6FHPq+46IfuqgQSY
kPQKOKwCzsR9GW5JyoXnCA6nqIxJfCv7EFyveaoJ//RUC6Q05NByLOjTxMTFMUQMfN1wN8X8VAgm
sfaWU8WrTTVzcihxLxpXluqB5NE3IesGmX5HkKs4RA91awo4RPJwbA43cWHg5lwI/RaqCX5q8Ltx
4edfEbspqOxox+vaBlqMQeXRlxQ6eS3zwmf2wQBTgAOWZl2ZJ+vCvbz3PC++1IDSfrsVCMSB60JR
g0gNkX7XNj5izvGbPSn3Ug0998VijawzYPA9eFyaP5BKjiPGd0AmX+7URYfFc1Z00uJj2tFYex5z
OhMDERyorMiyhOUq/Tf5TcfL2mCK7cqF9GzVFEX7FUEo71158zaTDmhpiLB7qS2WpB/0O77YVVNP
iygX7v5XRfIhEKlG/CkrzZgB+Z7cxQTOKizbQLP7DQilXFvFY0otyVyjMZHp1S3U476kBCCS3bXT
wJgfx1S0Nd5TaRsmzmW+A+cDJGj4FYpg+pfF14ybTtqavpEHFkQnIWjvn9WwZk/wRbLwSb3O25em
bM2rlwn2/vB5JtgVtcyNLCAWvXLtBFfgESIzVAjdAV+DUgzvG0zDGnPSRU7ZARqlSQaeeWCfs1Z9
rAamII2AFxp6LVFjU6s9g1GJT2bbXImbIC0eCENREJa3O9LJPQ8UQYXayg51mHlU/kU5djJidDIb
dOp8mFC0piplpqyBNtEhxQmLhh+RuE0M9dogbfBLNP+d/FtokGFfUrjN/8er7elCapqE7z0SC0Lh
BNqudHEkWEByJ9lYHkTIIPmX2OK7eypC5TvFemzl4lCF/hfh1cS42VGB3veHFdEt2mTmhUIgAgPt
cnpMSpfb7us7haZr8KxnlWH8c4Pm+YxIjEBIHCepfE3INEwynhPOAutAlPKuSfypkdFFluzAoAe8
r4VVeSsTob7gxpytFBzMcWoGnD68xJdYrPypOavpiqHhSmUPJqYoIaqTCLoaON00wIdWGPTQH8Fh
mJFTUJdj6BAkinIpaogRIktyBVfILQIo9HRWqzmi6E9O5Kxaooek3RlIvNv8YHg2yEZsfdo62J6J
0nj0Dua8Ne5J4tXVJLCYLxK7Tt/BZsohTX9ngwX0LPKUfPHXFDhlZ+mEWq906QSwhAS2DmhjqsHY
skGya5zQoYf08KsKhsQoNlQyohDAXUDXZ89tUt41cFbZkTkAkxR4LI0mLCyh4Kx5KegCUXMp59rb
J6hRDbB3U9HQYBzRBgncTJTV8BJ2lAcWjMjK/+cczkTBrcsgZbsn4V/WF9Qy0pmYLrmBon17V6mC
AuB6KpkXNB4vsMIExXB9buVBdqVklJpSYu1PtRTuZ58Vha3A/C+T3tsj+6BvQcvbZDH2tkouhpEU
KXTaA5LuSpfGil1ABLNwzEc7uOtma3WFFkpnaUzP9XhprObATNZFt8Kvw4HZ4p8XKVTv6pQ4tLvK
d0N/C90FmOTc9HxmbAuLPMvX2+XaQyGdlz/dAFTzjgSi5ZMtlZNAzCrNIXHm95SkFK5yxLVw3Hq3
CgJGABSSAEYB9MvDontNq1prru6h0LFAJ3tAkf794vQcY5w47NAxldMTIML39eCfqyCcH+ghX06E
413B1+eg3unc3JoFnc+xHWhSXzhOTshTh+l/hlqMzfU6ld7ILm19xGk3uPFBnM+mkIlaBLQGsGB6
clF2J+PLJ2wTe6J60QGTOlYWVQVGb0DYsn4HD/0yy4m6YKqLAIBvj/6owsuJriHJhPeW6F+Lteov
edvHKTZhbxPPGXI+pRBZaB40aUJqu0aRLLkmXWLbovIpE6nSL4oCZ+BU2VCKrWB4cch8TClUeZsI
ahSPgmx/J5PQVh3A0xv8SB872p0azuyQIDqHkw90kmxXHPWLvJ23e+3QmBc+C7RdL2CsFNYCZ6VM
k2l9jSBne0lDkMxu+llmJKyvtNR/M/rpFTVXdCA46OYC3MK0sqZxznwLOp03ZkjSkbCmBubBjecK
758VOKmqwn3NjAi/w+u8gKFzUVCYksSEYAEBZjtIgpISfD4t+jQr/BvF+AycbfBx/0TCughChjgC
DxW6L0GZbdDJCs0jQgsS7xC/UicX40UlzUh2pm/vuC35o/YO+6qwmDOsh7tnwbb8TXzADWsA4opQ
t2FrG1e+rgRmpzIrw1KrPQP7h5TjWmbccCtVC4MGudCjk4FoumJw3InMPTXpmkVNd38lRGROT1qp
A0KBIxErVXfAmdP2VJ9zzlc91cJ6z01AhxGwudR9Jp69y4imuOx+pQVUOkRfeCL4p77wEwq5zveR
vkiWcdDgBLD8Kmgm9loBdAEwrW2GoEzG7p9ynAM1LI6V4RHq2NMeOaixNyoiodlSRiMCaF1WS0zT
FCmpmu7LB5aUv0kn/U1gaTKP2ufNXBh3MugI0a0bA51EqdaP9u6WBlAcHk2tw+jnToNlFG2mQmbn
GvpKWok9Mcgjbxm1rTKRe8WYcvOYw+2FKJVUOtdTZJ91XaxXvHW1pNFj42Z7IUYidJ0CMAty5CIL
MVDP9WdqyQD0bxTJKryOdOC4mKbeCsse8WuKh6DVMZl/ayGaHCanN1J3jRfh59il/Ipu7OdvZ7nj
2+tYlLklILE4IlkFx/6deiaioESq09kNfSIS7A7odeuz+8HAUsqx4hEa43cd/nCrPxVgMxf1Brw3
hIuCjo9npIF2B6Kwf1zKmdKbU3ulrglynwM4hzEBcA5aaAGl99v7MWfmJyEUBi7gkLRXwdZ+0Ahr
kKFjpP1iploqFAvugvS8wttmrEStUBZV7W83J85SeOGZqRkW1IJ37qDLWWWgqCEQZgHyPIdSqVGv
BjIcmLV1piARzKaXl3SwyLgNNmFDo7iUpc/PiO6P8GhIEYgaNJnwUpvwXgkShXXgJ0f9lt3CurfP
JZDMFUwom48+4mR4nu3DIVByyEnthWqJfKsEivYD50im6AF23SYqkCegB7DOGG/qnE/IAD+kQMzQ
VJxjZWNeQag2ZyahGXNIvTEo0deaA1m7noBvhGZKJsXyF6QZ9Zywobcs+49fui55y5pHJFioPvun
afMKKPV7RxJ6q4D7weZoVFgYhS+w45ZNWFnqnIXY6wXshLzlM0JaXAfyn0lj3PBYBZ5lW56/FzuQ
TrSfX1ui08z6B1vVc8GHzCi+YHjhCZane7C4deL6BYGeyb7GGLvZaJHh5NKgSX+7fxhyAy9Pih6Z
9C62gYU15yvWRoa9WO8QVikLFOUXKNJpwVHEfR9VgD74sXfd3M4CRGOQ+2M8d7XYMT8/+FGL0O5k
mplUyvjSN4GBq36We/yRf3achxDE12K+pHgdTHbxqSVfHQSMOj68Zp5LP4JknKXcL0ntiilxoJmq
jDjPNYe0tjJiAMr0bnKzLk366CAUpX/uehdtLmRPtUEt1cgILGmxvP/f50Dq8rHBeFB4w7XN5yXT
p2tk5Hl6xaegmthpDzSxrhfyvhIHPwviBLlqNJcwKjtEwZBifxp8aQrj7wApG2d9Qek3Uvt1wdDX
vrD6Dc6KREwxJcAZ3ETextL7x/+NlVnx1X9wbVJ/dh+mgNZmLFzhCT3ereSGnzFTpalRhuXemoJ1
MysTDNbGXvATWkryI7bKt9MaE/EH/Bx19DubghfVfSgjk5pe0fJjf+cXwOIrafDxazzfF3k69gku
RzyVqCy34Cd6Ba2P2+VzXYS2//P/GhPvGwEP02sbGRCY5aOvGTCLA/dcnpVvPV+TmSRQ0RhNCS3C
/vVCnSFM2NZANDI9IV/5E2s8f9J9H572P++KdfG6mlVCB+DTeHWP3+Y8t94xHRrtJupC98xOxrvz
yJHNoR2zf5SNotFMWJ/9rbyr7UR8LwV8sjRLrl/PEfnhxQJzzIkAHURQwGWNqR5xD+2U5LWxpE8H
9vIkTOEdxzhsqAp+1zmF3T/eYfGw2Qz8F2royoTt+H/Q4nzQzsS9akmkwtR6dl0mLpuUN5x8IxFt
tNiPRjx2uXIUocNvuZfDMokJ5It8nzhtBJQbE9xnS+IAAtBktBJtec2gIVKiqkHjjagiF1J+cpxZ
elY/wyhrY+rbfGDHTauG9dbSGYosZUsRhKQcCn0ajS0bxZXeSsG177HpJJHYU/71KgkXuEABbCy6
NQ/ob+fVWVMne74T+XcS5gtuzYvOmMbwst4PgNvu1qQ1QrYDTJswc2zYnHs29mPTbmGeiHHuMFSG
qqJsfuVpRIcOdGKUFTRcbXXpgiwuLI/KxMurRdbtdF29e5wQHPCEVHc0kfi+ZcQ9ADH6zLQXJia9
ORJpHFxdxMTOlwYVKsyKGKvzwvZNifCBHp8St5YLPrC+Ob0oC9V7vVPX5RkWUM4k4ZwRvxVSFXRa
ZXxkEQREMRyUDveeKfPa/AMfdMTuLudB4FD86q/gDzQdQ9Tw4fCEMwmA6Bnw6jsabtW1nqOgMFLZ
b70SdBtOAQb5QM/RVtWPBOQN/sSsISKvnX/oaEIHuc8XUcyammpSA8daaxrQNYmB+WgSHcqGA9fr
oYxVO3PM/oEmZMqQuLll0TiSbkdFlWp81lnax88bt02KnA2QyEydKjn8vLuB9ZEXnUctTKwfrLKr
klT8Y23IeLt9nwXZh8H6Q1FrnWhKjFyW6Tjwv9jJSfeSokSlCqdh9hz6563dtfySQ70aXO0ffhZj
EoNHX9bH3wdhoykm9bsaOxpoN+Zeqjqxhub5zZ+YuGS8c9/PjY8yK2N1cMyno0aKQWOe8ngfZxtk
V7DYP9LJ7t4ZRISBlY1CAQQ+InRyJyowsixGeEQFjRlpFLdjSZ7F742HRAsUp4J8CfKmYKcN192X
0WQ4MabZsLZGVIHQnHT0E6fZ3zq8LVFgfIDlsjgXgbwhpqTVT8Sh0uCOWc85eaErqs1Ih5u5l/Fo
nzOV/QqdSVBTtN9mAq+qcaN+dc1NP7LDiFezpj0YNXbogXJqrb8bjvdzxMQngfM3ggG3iVh+O/Ao
9rldhQ+rDK3X5DUsHsto6quyhhYLa6WIb8Ot7v0i3ww5S3kpEXjPVA1JZdyTzbXYJqIQI1a402kK
Kgb65NLNwDoW+tsm8psNnnHfCR9ULusn7QCP2aEv2NaVWjImAHviEloNuITTpAxOYV8xhIqxF9Cl
U+NSB8tk8XDC++qXS7AqVqQmlCUrVCKE947Eo7ppJV30qBUASqoW5mvqVP2r7pbD1p8yAJd4oxaT
kMMJonYT9UeAqD1/Ll2AdcMbV9/YsXqrCqHGWA6rx03mMCaOv3Paa4m/jr+H/lNEUzHLtcfl2kFc
Y1fA6aDNaobmXvwZlKaRUqj4hUoUBEVzF7Ecq8h2Z7r/4qbPftzP+2wZuqXLQEjLq4CUeZ7N84jr
fZZqwhiv6egnc7tb15SoFP3QZlD/R7nECCT7W8pGo9MfyYmUDpV6WvLWiHXvMFVfp+b7EoDRsd4S
TG7eSm3EJfd87TLyqUzh6bVwmI54cMwmML48sgiFd+lBj/PhgLesdqCALs5Jk8979U/6ADcTbC3b
pkS/KenYotV7D/LIdGLFqD7AHIZj6gyeWF41ttQo++YWkDdGE5O95guEetGhvB5ZjUvDIPFi7/KT
xi664bG0Jz9dyGAAKC5Qh/omAtK3OQASNeSTGNYLmPZInipgJIVrsodD5ZKG2u4pSnFiQOv7SIpA
PgWXoK4GHBgW6sIwc94Py1pITwfG+cReZPmgZczjGdd2OqU/4srAxX6jOwB+iSo9fmZyWdPQ52mj
eSCq9uDloUQPJWhULD2oFNd/ZjKkDFNRe0AY8EW3na6nUK5eqFDGzdGYhh1rrIqZHJdtVoh0rZPm
G+Mio6ZESBYY3/15ZiNWfaBPJM7gt1cnN5mQF0iP763lg/ITii3GrMYL9WNN80xxVzdijo/utJgQ
xYxC6hwFiC/Diw9C9LXEqolvcvqlHHkwiK4nZJx0Nm72T6/2Km31xMKnXMi04riOk67+0D9Ym9Va
wV+kYBpfcYrGSF7vUaHWKGwnm8jwa6IvwwLNuo7h588mzssVnTzJ5GuhWqfCILTqjHYbpFrIwFPi
kBzv+jsFcDDd06ya7cU38YNXoC7Y47PqBaa0bfpBt983iSP4SulXWMl0lewcVpQKLa6KsMdQMQ+y
fFjMmITIjjhd6WFlsAHJT2TIK2xi7V+O6P406F+/y19Zv9gzejZNXbuHoAUFdx03mYnfS2l4oOC+
PqI4icdY++eH3I3mxzK+PlYdn9lFmKsWIHJDwlgcZan8E4O6NFPptUWnSVlNfHQLqo7BQLFfhBtI
Urfas8wKufp7xm8P1mqdb+FkteXrRJdOSYrYzVrS4SN2FNAw1JHt+SH36Z3QaclUTKQLwZyYKfzS
EypUovfiI07WoAIh4ZtPuqHjuhhaqiFP/fEtxkmHUd8w1HIF/5gQMgBVy2G4YNU2JbDJVSWsn+X5
nn/S5Bin5At8tfMwgSaTHDNmRh087jZnD0KKY9y4vOGkSQPS3BpNe65xx4PSDYr6n6gT2WS/hp6X
NnZEojLheqqSszgZ6pOqDeHKgRny6A5UDZcyRdhVeDZ2PuEKb9BdUAdA0+nc61RegSsxsPYhM+eK
T2Di1ZoVbI/HyNx1y/y5CaEos8KZ+nxz57G+rygot5/ft6Uv7gzWMcBJzCOoPYByZCdCp60BJ0Gd
MZud83sWDO5r7/zp9iYnC+LLHm9I/peFfr2nmh6+H1gEkvKoH0trSD1rl9XJ9LzPU+9WyJ1Ku7en
FfFd1FQ7AvAAPCQZ6QrsIrCgCcZD4CZ3Yzl04DxJ7TVWGg3bM4PCeubuHGrTIOU7Gkw5ahOrNo8j
2b04lewsdqwJw/YTxuejkVA5lWpbNyD1LBhmywYFoz82Xt20VVaoGN5qPDNvj4+oHiiGthbcm3aL
if/oTxHVvU/vrUhaaQUaSzLY6UL7uf8luh5m8cbDUH87x7+0w5pCuOdULWfHG8/2Y6xnQTkfPVQ4
e273XUdLwqtq+aKgTK0nyNok9V7C0YkSbej1FawXJeG25KOzM8sKnuf7X9ZnupsKK7fE9EYFqcsN
cW6EPLHG2BGhLWeo3MzDWqlQC8AuUupxK1+MM9GUhMG8EJNd7WxEqOpsNi+bgDzLJgiVqqtAMmIW
hj1DdYvwsgqQt+9AWNi1qH8MzuSCQIKN5STU6FPmM0mDzILnS5q1BelO4YeSROTLI3bmdtcQ+mBi
pmTNR78VFCwyzj9IbBH0P78KaId/00lWYEuRq61H0ai+bdrjpo6++taGumV2iGG+7EDRvrYU0chg
Gr76xnQmp2xdeFLaLoRE/ZgraIEEyoi/6RE6zECE0A7ORYtVPeefCzD3PEctVcfgzVdUsDkuJsqs
yHVM5L2hoxjus+t0/HlEHq+5TzTDgcCfc1336MQCM3Zu6KKgcwms3BBBjnLKRymJTVFY4xWtrCTO
Mg6aP7gzU7jo3QZUMWE4iWeMlgvVRQqwQMz1Y2Nu2q6udomrnkVhTPGouiR98HuPdepVRtx4gZfT
M/zi04Q6Z0qfCtuRmAQ0sLM+SdjOVEe5cRSVHM7qaPwoar9rfViWXYV4lg9aKs7VW1Ic3wTrw4bn
a0JRwqJ+zlp9d1PhUO1WHPjTQcLh9y//dZgJDCiNqh0jh4WAqWWZ5YaDGBleoT4LGE3wC+hK/DkU
yAKqz/viJWmpsqkkr2aK92egNiZpOShMUVo0X1LKtavXxFMYC40bc4Y1WFzIzLGm5k5+JuQv7NEi
lLPNyUy/8UktxPkJyXkjTGJ48EhAEvdzh2174BEUG2j7vOfT4zOnwa1xFy57DtML3F+8I/oxN0Sr
UInT5Xn7r60zMOC6Rp5srfmf1UyO33LB+a0pR0Hd23uc++XHnj98f1u9CMYGrCTWHbw0NZXChv/X
uIPPyhrqK5zRkSqGmg59XdgCyJo5kPdzzb70511Hz4mCMiUmAhPOcZCxFQC4aEszkKdOeyKFhkOv
leJEgjq9+aL8jah/BCouYQkyHbyEPmaBZihZNVFvHqKPn3Qy25jLhBi0td9qz8DdmyKKox+V6h2d
HRWoS80wzoWs57VzvJn45NGT42kjyfR23Bz421rz7kRmZEmfwMojv7MrGMSXZbZFsuIbJKjhXlMD
N1fGLA/WzKOdUXRoaQLa4pdYZJKL0E75fve85M3gkf1w23318UyHCDxVYuqD3K3atA5MazRg9R4b
wcmp7gGGGH++rwXDhmWLnP+9cphmwkMgsrP869rk4EDsIWWoL4tKaGllzvwP2YDpjgjfFenBBA30
To4mQbPLsbb9NyXg8h1O2v/H6/8+eb+wsdheVtGG6b7gjC0YXxl/S1BHnvfGFb+Y2XlYK31CKXza
Ns22Cok9zleMOETQ36xUFKvfTJ8smwvaNPiUfFXjxDSpWYIh0Gray4OyO4wMFAfgml2RljIg7XEG
RZI6BLuOwT81BLnd080eq6IS4an42TsFRMnOFT/+3rdObTSKjzg0SO/cjtOdWYCSpma/mf4Oglj1
TSY437W+8EsLhELSdkyu1El+cn1nun0Wh+UobpDFynDrFkzXIG5CRtAFTd4mo6WdHdbXouUK+6Xv
ffbQVrfsiGEMpxpHnEgSjNlA9qINFxTOgDoq0MLqQx42zITyP/8gEaRSolH0CQ1aq2u4eAzkXTtv
Dr5I4uJeSjXulJ5/oV6Sl+3Hv5jFYe6+Xw8rQHPKr3kbSBoIC6XF8FvkbJI5weig3Yq0HR0CYhPe
RMGK3d7/5DmoKOf9Y87B3A33BC7nMdRVVetUqODv3WEvOdfzCr9quXEkQcV0ALJZgmdT921xybGv
3xD38/khjbZivXxENv5sxaDSd59c/2IuOMDpB5Zwne6iqO1Xbqw8a4XnOa4EKS/EB5lupFfoP8Uk
85X1DcQ1NwFgNXmWJ2tyGuYzq3OE67fysDVFPEB7YF6xDhoLUZgLssuglBoixMbLsiXb7f6p7r2E
clVVUWjBQLyfzJkWTi19hAs5nIWgNv6u0OjpMVMV0Vq+z9y6UmRPem3dHdoDuq2ZsKkKdDgDcFsM
RRem2xxoun6CpfkTn8KXPCOJKgXIVQV+EXYxwAhq4Ko25+bgm19BZ0CjCiKKfKc6ISd4WljgWqnI
s2bDOpw1yyzeN4QZ/qzu+BeBs0QpAgAVgHjhSXM0/ITb+9sTJ5risDq4ublaGELAOFb6M5H5DrAl
/uK8iaZzk/f1YTljg1vBC9kWGd8V3ugFNFiBAdOc1ROIFvO+t54aAGesNLrPTMemNmPXRs/IBgIp
rH1hbgptTqh8KMe89ZY8aCBbA3jLLQJUaSx9VH7dI59ZiWC17IxvzKcJ7yORYe+YABSKuuCzo5iD
j+ivYiga//vDphg1rIjsm5g1r5/dlsJe5RIjDbBvifejPDkZBBEX3rBOTULIuNOO4eBxtqG2d8fm
5v+1vbJ3y7ibFtkOJUS/BJx7k087tulvI3b2aGscj6a8YexhbKtNUCn3NCSkZYRzatufqOyJaRlH
bagSF+dRYx6fINvIlAZtcvjwdf/YoW0ioluPmxej/DqU76kLD4xzf8qmCg4ld7XYC/HSesK3BTqW
6+Kp/fg70vZlvmhP7TBX5wIZwdmFcfNuR+2Tc77V5nC3+a/v+tFJlTdbaWRz5K6nX+jR/mNXSpc6
lblPF7TEDqL65NRpdQ4hoXOOHc8OUYNKh3zzgXPCtXiOMkjoxSjTXzVmaqIuLpx4M9kgHFaHrjF4
WcV3SHZD17B8pM3lR2k00CSwm2w24BG5JhMu1CnIB9pfwdeTxAt/oWWTZc3DrGd0gV7K2idC6adm
faHGplVp7iHvFr8+NZ1LxhoJnBz8cy+Uezn0Ehab82Gk+r+mwFepbjxvq5rT/qYuDhSjX7n0LojZ
oHR0dhPsjmNkcN2AvjzKMl5HPizuV3Mgu2FvhzgOneq6dnuqeHTAzVTDvKOZKKJ2+/dZPK8priHb
xYrsQPsSmpLG/2iv9cCDwfLkoThoN3U53QXBsmqetdEUYKaoQJN0ZPd+nwARzSB/sy6gut72ROVu
Vwi9g15u0PjVwWnOxvdCKzfBbQa2MJ7Xjx/vJsnktm1l3DiJ3L2j2+uchRQZeMHvuSXpZinGEhDp
aFVOZ4nMAByXgqLKW0O7RUZ3YBph/70ZIyJoad/CZeZ0XFe/e23O2V0luKytEBFyBsG6Gjk1AZff
FJ7KdL7aGoBFZ04Q81ouPAFfHerV0s4E8AIQEKrkbQRBGOzYBR5IpXf8Pi1Iek0PFoSsOSOnMo/a
rvf1Ddry2CyjBUThaFx/Pe1Vl7RNxuSTCNbiSnUR43axBgB1e/i8m3DpieDEoKRxvGo45gwzEKw1
A0sZW2ZdKnCdj4XRMy7aO7H0Yhg+O+YOAs9Q/5HjHpHTi93VeU9TBg3UrOAGecP2Md0bKVrrnNTy
yd/xNzT1wwLc0YqO0/n55PgIkqnMfjDW27rGQWMrMDpLsdKk+I0pq4DEt++n52AZPVUSOtkxHSlE
2rR3Mhv3yDSK7/fCyGci3eu3Aka/G36mQAUlj5DC70xakUoEAxYiwDCb+Gk/Wrwuzr3dtSWH/Gct
r6SKMUWxB7TMzXtRpx6AwhClcAt4YM/R9nI5frhS1OBAt+z80kI8dre6GhIIS35g30jcSu2Sb5mw
ivFY+KQxQIMK91T9RS7GcSquPT5ObbhoIJLMxxhj7f5azC9gC5zYshwFh1xbIOmI/DNLL89AMvWQ
TvS2xvZi17c/e4ns9ZyNCLUd8nPw2JMiOQnPq9ez345W8EYUQOHoWHK31M9agI/160u/gF3Xm7YM
EbPGG4a7GNANBz8Aah6UG+es0qQzWpIMwpVFVrMZGxMOuGhn/SQCGWj2lKUETc+v7bT9XzRkJAsR
uyG7jYSZD+Bn1Qa/8fNl6nXr2qspBFCBpAycDbVuFbgw3i5e3KiN9yH0bWHYa0IZLLrTXHcZ0VRR
pFUNiVNPeB6czznsER/EM6KG3eV4jBQIUXsJTTcx0smdLTXAZAo/8IltWwnBo+6P5Sfys4lqgeWC
Kef0FX5NbhVfUyLcdNqjH6elKNsJcbHPgi4KygW44v2Svl8EgeJ3Wrgx0KSuAMGTfU4cQzobdbUn
YnEC9UyOc1BwkHwKUb57UVQf59G3/fFfFwE5qPl6KDtVGyC+nIbpBxMaNvzJdmeEBc7XXcdqpi0z
gjBsq20A+7QGTQ9wUjjQc7KjaVu7pn7wvc8UQZzYesoGMkKMMotALsI8dG2IDR1CA2aSSaqHWdqf
KiEMxXL7VDJn1HH5LFXhXAfIBC1EAYSmq4A0Ie76iyJPTtV/hCFe9AB6C+fZJCU5Fd8aBQJSim1G
ZXydQqHKHztho8oAQes02w1tK1t6PvZXIS9pAq9OpVKeDZsQOveezaIA/GYansYRN3PIe4dulHUz
jVNHulNDdH6gocyeNtCS2vW9QLiaMO3+GneU4oHO7uPAlJS2PNzMMXOfExU/WS5d1UgNqehBHEK6
EfKMjhh7HMmp1l8BwiYtvruTLUs1Jjg6fGKVzlnRff5w/H4R1G/PceH/8BqVwo0jM4AqBAXcmgTH
lRcWeRfLMkB/Vw0ow9jMR8GunPgVFSlus0y/EzPMfhCuT5qppij/SeKDcdrU11MIWLyY6/aksA7A
vN3FtgdINPVw1M2eemg9CoFgPpSE7GGF3to4t6LH+vTJ0+YpEepx9iPuRFUyF+uv2v1/rS+sT7/D
vfTWY7gVndvJsap3X3dv1EicAWi/ublBeJoIIcNlInLdp3US0t3tedN/BEvBnMzkM1WOuULxrirr
G0SsVIf3y2JaBkDz5nzvf4vsKpDWbk1C3IW5HyExLCJ1kaWhY0lY7Gh6N/bv/vhRuwfloNg56uzE
K1DtTpVEU9jOY9+G83sJ+Sbqnss8pgtcweywbMSFkqHuCelmClNZS89urRaP+jdNQQbBPjdm9Yw+
kWjh3BUVc5xytrUQYxQHesBLq1XA3d6lsJ9JRm3YjSi0twzEyK3DxWJgJaefi2lUXlzK676iY/pP
r6Ag+Y9w+C5NrzvnM2vLSrymaQgr+cnsWKr6kpOIfrMyAjGCsxpnet8l3cBYek9GcLe3d9Kb43NG
PzILdcoMUa8Ak1ckxKFwQsbSTVxo0QZnKY+135YF1pxiU7UyPxujXzfS9+K5k5LlFVPPdLKTUG60
gOqW0Nk6lrIKr6qbRLq95va63FoKMxMncha5wqaGj+kVTFZ5TIM+nSc9BvdPUt/kuQ9tvBgzZFLV
TwT/f9+qeabBpyLbJ5Sj9yhgaPriszcQTpakrztHxz1pJjxDZVAPfym/NfAoj3AEAiIyPsWLsfPl
Xy2VRtjjZ4nZlrh9GGdHO6mXKRKTailYew3QUR4EBvJ0cydWDIxpojtRgPKnUsE4+gsCMdTD87eh
hCtkXD7U92xLNafe9GWDoxW/HPrSjCy/NfgWx5TpaLmUof37S4RR3uAFRmY4Pd5dOYlUc/g5YmXP
mBdCUIOZFJ/qsraU12QBlf3x/DZrgMykKffh8rNal4qo0qq54NSpemt1NzyFWwFBTcUDkJ9UnhKU
R9aiMV09g9ncGrWW/Vf1kx+tjBleVxcfqwCucm+cWD5Vj05OODmlmLR8Iiuod2qPOuNHNIB985Cb
bMc+fbMQPKmocZxnBVoPgBfDUEUoa1PZyGk2CdOzLP1sI9pPjK9ABLBUWk7n0tnF5Rp4sLK9Fhtu
Z0lDCx56AgvtgSD5ywEAGs8gOBco6e0b/HAdCWOHNeqYIc+Q/s6+0FolpBpneM7Wt69wPU2IOWA6
PKZwC85ri5XYD9SQMw5Y/iB3nYHRj/qS2iO2F6ZXreTsSaqwAfdV6nzx2+MBDnpHNVOo0Jp6RGkB
ML+5VavGzQtoxzNzCdg8jvWJGr2aZO0h/WehX5V7ZqmeuAmqv4dzGTXc3Bm3S6Ulndo792CRPopF
rsZtOxVYPk/QO4xRgJCj9P60sHK8fR/Z8nG2AiXDF/ZqcEoCEeSl7Kol9wZZ9O/gO2G+9kR0ZWCT
OhlpByB5YJtXuode0R2rMI+IV0vEhfWCBd3ukHycC7GyoputriEQzsEK6BD9c8gzyYf6YNcrMF8K
5GxVaTuy2Yq+F7AG+/JMKUou6sbaKnOrnZ44ha99qgvdWyEYnmD2QU11poQYeXjggyBeORze0X35
pW5T/2NmBgdNfUlJGjXZlt1MxhW6j2hTr3GMFiBN/ON0fpUm6haaiss+/vhyoXqdxRvAT7o/iG/x
m0aFDQbQtp5cfd1GyA6v2U+wDX3XN2576f8EHQxwMTzejZPTsi/cFzcUTw9hm4w2s2lg/qCEJfGv
S4I/NgDRlvOR+JyPm0S+UbyyDWLF3E9YGuPahDKo/WhyL5HEOfa/5sW/pOTyWongbYefGEP6NwgJ
GHPxIe4TYKVGaAA28CYzmvI0Q6Kpz82GnU86aSGHXIc4X6ervR5tNU5wkGEWFA7kQUut6FTb/vUC
wz6a1fIkQfj29H2mqc68hIZKfG/foc+PpW5a3QvD4wKYVlzv8dbxXJ8WJP9YoBw3l3e/2Gfm6MEJ
hbbvIaA6mmuf0uOvh4Xh19oGvV7Fox/yqimlqVU3zWrRdlCFz5hC0DjdKLCrDuu5STXy6d4niqTY
Lo9vlOMK2AZfYDo1g6tJZhHQw9VwlECUx5871dR7YY5gNpdIFfh93YuDxhqkFcpnPh5kmcHG2A+u
RMgr318QNDsp6yyTNlGFGDvCFZiZETQDb9IK2d9m3VHCMA/Yq1KmuIBL7z2ktDx8U+ikrwux5Xfv
TzbftxiCih2JGhUrcQt/fRkHyII4m4leexhTGfnCAtBoq/v7BDFAL023S6kn1Tw45Cyqz1WFcSeF
s9tJ9x58P+IQJdtpTMJl617JpZw64p0vgbi8YKaDPTooMNp19MgLt3cUcn41qOKB1j7gIM6KwmYi
vNGhN4YxbjFmDI6XgD13mS5vh2zT2sFMu61A92hiURz1s/I1XEcMRK4+DUGZHAAMsg4REgmm1j5s
2aW9vVVO5O6ESN77Kz6Y/ZOrcqFfH190YIy4hrDlgMjqXk0aJUpKXJhhTXiEpkUcKmz8OwzaWFgh
j6JEHOeZW4u86GzPfQgzCRAXP4l9gEiWlBHjGJDe67FbI2HMO07QctOCJWu7obeiyYTbT45MuRAf
AHocfC/z1gMxwBfuV73oL7DoHtF9tzxpaqXl6M08j5r9TNKp/1DsXGOXNnV2yoUY8TwVzolaqpkQ
dcqMCpSUTSLw6aCW7Wib6lcPaAmpPzTLmJLJwfw7F412jn6L4ihMk1OGUmCHr8SxD5J82ttIOczQ
YpfBOoKpOBAK1lSAklK9pSHo+knmLvD8vxR/byajx8zjd0zPINR5VU+JNSpqsGtGNMMuqsz8yNcM
S6+tmLtNWabAymqdgeL+8Oq5o2JekyBu78crBOVzg0axBCenJEmB1jnPynio8DoIHhQ1sFf3iYmT
SHpoby+GNoxDj77gQjiaIY26RE8M6BIKtMBfvkRj/tuxbwn/+c+qYJJ6AgOq1zrpeZFrpTMPn9+S
ZWY306vTqD4AbsNW8zo/4MCzTGVlqArOHTuHUavyDl8fTmtBCaw1nLMJJ4vaIcCCE3cGs2acvCDE
QpWERQBIOu9lHavFrPLwANGmDih7frd/fiaH3B6M1N97Pa6HE0V6nZZykHiY6l1dVz5GyB9un45W
6yK84B+5QFgCWhMwuz0XECx6TJK6Ae7/6NE7jhgygO7gcqh7BlN0EV0+mrAD+Jdf9+lBx15jA3It
7Ky1dL2Xi8TfIA3nmON/BDhPszwUxlWXLq6sYQl1qdy7zelWvw5SYBo+/Ng/CwPiX2+Lyp713PrH
eFYzJv3kpb1759Lw75mdLG2usfmHHJejUy9dLOWBEK3ySlBwDuUs7ulGcp35ANiBvswCVPx5iKfw
mMtvJ4OEHHlaIgY2pWohbxACQVGSIlW+ifT0mcXOE7oosuxcda5FGp98daaDWjEx+UniKZnartTE
FVdWhE4GclxKalTBTvqGTXEbaEVfgu6BVuzc4krsDkfBxx5lTbAJjtYlyKTxR0q4KYZgVxRqg+Kk
bZkPRhjzBistpiiSNVefGJdm2p+Zn0RyeaT7BGMf9nSkov0Dc/+icFsXraWUWB1+Oq/5dofwzm0v
mYGLDoJAxXNcYJqiBwqMi4o4fBaXlYzq9nh8LnWkB83HtaeSpr+LcRX5wXuft/OUswyPsALWCDhH
iquG4tofrhbMLZ/3IYMdqvoqXIb/kfJlD7HIDK0TAV2UEh1pMirRtABVa13nQUtbsE41PTOXrw6o
VsMBN8xaAZsr6mb0UYjtRdm7X16VxKGp88dvsWc6Zldh8h27+dchxhg7liwWTmrz+UzGPMy8YjrQ
XpwGN6nDNBTCKwJjviRzW2NH+46AEUR1d+L8UYvfiwCX+z7BQ+KPbLnBduCeLykO3Su+OsPK6D4r
eqKAMIIgYiLgD5cInICvtz5AqJ1x/07pT4e/rT7xHajjatD1a99s/+BtaSI26kipMV0EcuVg4FvW
40HAnjYwFHeidaZhgQbVE8zMuBUtH3f41jS/Q5mx/alfs6B50dg/874BvvXTciUKlxN5362BHojO
7sgs21bb/pl19xZ9uTON7MOItZ6tNDr3S6kHdm2Bw6dVe0QxYhn8RTYGTZulvjgTO/nVl6/BDIFs
R/N18Bsl/Tc+Mu0SWG+piYkblY30sOwT4OsEyvAW8Vck4UMhjaoZoz90iQ9tuHrvrohS5lGCf4Cu
bqZfC7M7wFreTWtnEQrGpGQ+1+bfwI/w+DIMEQnLuNbp8uwYdbBpyirfIB393zxolEd72n5I+tie
+jSdBqCneeHDcUYFxR7ZU2ugpWzAnrGg4N+8Z7Xr8uAbUQGHKQiZmBGxzgGVXjjUoRY8YS9DCG1t
zWz8eYSOyV3akJPkDfHGfjD+djE7ljPr/xxxJPIyj2169vy1RQqHnEG5ETCg4gx5k8Cdicdr9G7f
HQP9d+NrVcOuCkZh2B9dcZ62LcemhzoGmz/dX57uHHgbhNXEgSKkkZ+7WzWAe/1H3M+9GBvlPwRT
h5lMQ1RwSdMQL9WXZZDCHmIk9SOYjj24uZef5Qj4VWkJtuJ5g0Y671jvWu5cZAlL/YQk84kI3Sva
1NlCCJ8+FA1+gzCxMqptWGrg2CezfFBYsyz1ad+epf0zfwmCSKzprSB+h5WEW8Op5c2Yq78CdwTi
2N5o9wv+UKNa2bVgsttyddzveVGWwcpZKTFMEE5pS1aML/bJd4mDqy4Rzw+dqlUnbiIJjfz36yfw
mUfdKrqGP0haAAUkpvYE3+Eu1MAsfYxKqsx9Y8Wf0Ig8JLlvDwEE4df/YB2Sja86doTTaJmYlxD9
uq3QBNd0AxjaQxalfYNkkrH2/yM63nDY3X8nRijSKnav7UURmTp/RlwDKD21hOhOVN8d3bGeixdV
MvwKPleK32Wi6+FzqOnc92XrP3qq1NhX/awzK3Q1NW0lVxZoqLH5PWsRXhbu2dJbFM9T75YJxmIh
+fDe7I50irzWoKeLnSOABy7m49I1a4HjB7K+0VJWQ35g561XPwtloMlGP1cAzodYpycN1VqqO7tl
nnzzrDWig8UEnMW1M+EJqUblT4MDivdaXHafoxYNpAFtk8Y3wTbxASKLKyC4Py0nbgbzla7bXmQL
tox+IXZ+byO8DXq8eJGYLpjkhp9plhLGa2VOhACi64NLmz8z6vxGeyLu4OidhIzmgec7OaT/onPB
a1/IvTL1DsBfDNAsjdgjPCvC+ZknMUpq0/C94xN8BILpkMU/IKk7y3U1Tk3Qpng326tC/1EyrtW2
PdPozOIXww9FwhymP85D/zQAUHAYfRFgLV4WNlExz1xhRtIJjFzkSimENZGR/USzYPGCar9cAd90
pul/Xaxl/LDQ4S4GDHXiFJg6Od/PbFLL+AiV8lPCRPFCu2pWWlceHZtsvI/MEVdSr/sel/sJ89cO
7ytKPlmTcu0D7x4d7arxarOOezFnhrvO4xOJFirYuNMTYotPRrY+RxIcjqIXJgNClv4cfb8vsYUc
EGbUbU8y7QrDcIVfEfmIRF9iKlBNP7jbU3zGKpcwUDGgivlj/TkKiPBmPUxooEkoF1KQ8qVR2thR
3PdItQQu98ky3LWrpTD0U+7HppMz8UnUa/e4q4AzHBX1H4xG5AeGwfv6OoTLARFBqnOsP5fC9bVk
Zk8aUeUMXDYSyBPSs779t0ACD3+nWY5gw/M9WclwUqsOdiGa9O5Tcs1jHgdPrxx7BPzZYQeaIIgP
VUaUazIjCJUr9FVVDuvyHp3M38/V099yitj9QX0QYJNuLNlQX0lZg4JHoMw/A0LYayawUXEPVDfE
2f9Fdv9mzuhwSSEh9/hFUIKmjth08Sl8j1lqns4n6hDZjFZJpJKM2l8IpafAN+5UOb3Bqzh1rks9
8g4Eqs2izGiYbxfgL3goup13coWTNmA+isJcPT+o+Xz0PTfd163WIlxWL/p+F80Bz7V5L4PWxTXo
19ZRqjzHBMd3L0XnhMaopLH04K8o2Fuwwd/kdsrjXz7lyOQOAFPeMcq7lHqYI/7i5ZPLioJi6KSM
WAks+3tXTjooUzzEPYrb43OQ4YU/18fQvEjo20aeEw/bLrfI02ljckE6oNl4Djczv5tDDZXiqKi4
jCWfC/puQIajdsYLzNxMUfdgi0BZO8BqY/OxLiF0wU87yjtpqivK53aJNNHgGsOb0jgYaT31pjBg
Bk1rDm47lI3H1MXzQ6NsVlBy7OS0HaUfN2EcFmsnlrn4UrdsPbWgMQvgcsbqkEuPLebZTEL3+Zum
vOJT/sdHxvnUpxHZvYuvnH9ad4KQAGwPkdbmAF7OOisUllFXxJitikEhjK2ama7r326wFkbNG6ji
UUJueN4OXua09QnviV6ku4HyT4H4rgz1b7/LAYQmZ0RyvLz2UQq3jtUU5ZaDdDCultWZzRAaNE+Z
eFZq8CsjPQhNOGcWTj71No8WWfAAZyeLnwNOuR6bCn5Wa7FQgLtWaWwAHMS88uIBwusyJGlKXFgj
koFVG/A2e751UmftmskYGVGKJdE9WXhxMJ+bOjRw/bfDE/RChBhpoqBr29XT6icyo9o9mbJKkV4N
lJ1sGcqBpqkearVy96fQJHbDRJGyqJlmi8DEjFDLjJ13HfpubacSSo141avFpv/SopMpKMbGH1NR
RB5+x5O9Mm85T4q4XHwxhBUHgvsFxyWKdgEmVVXRatGx9DJS1GIvCrUpf6gsc/lGfTv6sNgA3qZ3
c1Ik3XrveQScPrmC65PHmE/hd/QM5w8rczBrKl5jPzxOoctKDzzsKf9Uud1zm+F1bmMfZ7FQjlyx
cQbzzs6zvmYvqTQZGotr5ZX2cKnQp4CH8v+p2BPw4HWgxUICE4CF8y6rebDm+IZ8CODq2KLhsIgl
/ICUefmJjzDcGU01IYlyhk7O0bP++E1kqIRCR1zjXvob4q5kcxMGajLH4bxKzuoS6u0BwnX5yoIG
sGVBLZ/b9UIQItA+K1ReybPqDcR2uZXOwsM43x03MSvQU7HtBwdC2ET1EPkGIgjeXtI+NC7z0N2v
mdZdY2O6QTU5h1dZcKAkwjZDIMKpGUzZFD6Zat0JvkCs7ZmBaWb3eBnvRY1E6XOBorxYQEvRoi67
BiAZS5jB+VcqCNVEuwH1WzLg2+Dmzo7/eDu/a13XROawtRWMerRyddJoZ+tdv9ZO41f4gn3q1dNk
UKMQpZ2VfUhnX0/ZHH5wD019Blpj9d6hGcHGefvHSrg+HvTM5nYhISMn30bmv+2nVT3S+14PQ7Yk
M7s4fmuCB+rWTbSDQbvv8k6eEXDBh2rJ2H+dPjef9gnKzp45MfbOXZk/s6N072mBssNk3y4UrEoh
HJPmEdl4FQVT8b9TdBvnFv03eaJSsWz0WSJRg2+xEqPHy77MbJHlUBSCTB+ZKeFK61vsDsCUTHlH
dxBQyb5Q31/oPOz2GRwjwTc+g+VefS3lQK2F+TXtlMf3fW5V+zih8D8UrlYfx5J2pi49ih5vfa2J
RhTlMCIvcNLNEw+q0V9REZpFUqa9X6lqTYBHluLP0He5O92x8865tPlLt6SDKLx8//hmxBhgEBxi
/mILigD1pYKscXIfACHyCqGAnVDtd1YkaocvTbcx7vlz2SvxDrvPTXqfxK6Dk3VYhY1GKIy6TSr4
yzP0ijJXhTP3nnLbmujJO4MBMg5PNuZHWd6SdeH8foJwHhuHHt92HpOKetO3+EnY5ySA4pdQ96vd
uRoL/nO0u+Yv/Ul770IhwGedpv5uX/Nt8jutLj/k5IPuOkP4dtXCJ/hwAIkciz2FMkkVb+zV0juS
vBsmtAmrhS7ujOCG4hvg5TtYmoMZRt0SQf/C3/3rGUWs6lkVJIOqYPwbVtacdyPrsRacAkzAMKA4
yHnJE0il5yXEfVEitJi9BXkFrGrejh0Zkmgg1eexkjXj/Fc1iY6/5o2jGOiCE3JCtS4Z01+z+S7W
PImPZ/XiJlXK60Whv+C0MT0EVmP90HYB4jcv6Ce6heeyIGY7xQy79IJqYYQcKQjIK45en9wQ6lCZ
K0zsPA1BY01pB3rJJN8xkhtAzjEQcF+Km2r9GiDRgKOLVZvYHdz+SXbjHcUYKL2HW2+zaVFQnUU5
Udm/gxPmZ3MjfaI66vgLhB8P28U1qMOvRi9Icg0YSztI7rtzdZENGFaxCSS1HeXv6q6mwz2vz5SZ
gts81wV3Di1swcmIoGWn2K+7XoP1Xfslue39PIjzrRfnoY0CdtJnlQkcLfK0Et/OENi3K/GEFb8p
Wb9AXIcLzJWJP3SdrY1Qz0A7rnASz2XzTTh/NMyLJLm+78vDX5PvZLDMcaRmrtnsw4eRTm1fOhbz
qlciAZJ7JPADNwucgPd245/3EOH8eOr8ZBXylnRSxPDcbW53eRdkpvfz1pWIVVWok4wngWXXPSuT
axorUk/BexLDRhQgLRyZzn/dq42wZ7g70wSOmoPh6vfz+3aXpGCQzbpuzON0mJ3cG4c2O4rrSyH0
T7xl+MtotjvshMFucHKLK/iHKpjV3JHQOsCJRUqTPoC21pu0btsdazHNRtPm1eMcyd+MxBvuHBCW
VnLe+MQqvQSExCW2huOz6lI3FNYUBMVPtDPWS4Y7LvafFxb7lNlLpgfC8z7rgR5AWBjMPOpb3xQ9
00eZroLD9hBzvD2a8jebgVvu5nB7BBU+cRxqdylI0o3U8xCA0nAoNYVH7KpLL8+9cJaD4u3dnm+I
qAUE0xBCw+boIaP770MD40oZOervg/W+WDWG8SyBPwOHR3ESsI2FH5nMX33eR8BIMvr5BFSMxhjj
78y75WkMQMj5athzynuKVfQ++uA6AYOtRBgHxnzCz6ot42ZbmoQLCC0c3uot61LdSM8rSX7VoAOE
PsXp6ka0Xue7tui58z8OS1jqLz49vlKwzupmUE0bpq2oxEWJLIDNrfpjsqndFE3vJe2JFW4KDORU
6VlKF5RUCES50hiDB8pRTQPfm+JNO2vfxXG2W+tKtxWvg75skeIfTMoX/rV8nUZ5trT9l1me/mn/
sON+Ri+eilwHpd5VaxzXbaWrkq1BOlDACFDfF469BLSRpqr4sSaTlTzVypVULOO9U9ziI2nRHZrY
BIZVM9R9gjHSm33kr/K2ozcmgFFUG0ASbKxnJy9QLQGQnvy2zOc3fZRzD1OPbAQqnF5j3YlM4aS0
3ufIgOkAhPHy0t+zbh0WtkAXGs1F6xcv2KzxT8ysz0PHiT0tcVmRxZuMLVxKg55FSrbx4msGJ92G
coR9umj7eHgh+zUoOWcRdZWl4rSOALEqmhGqAsUJhoH3fXAx++uxiZTVQzANgaKF12OvnhjnFcJI
nHKomKFBFX26bSu08ZqNgbmkXUdwTDQNEQ+vW8CYxVR8yy99FCuyIQLYzmIiiCg06piBGAE2+5Fi
DRT18FiKIIpt8UANZfsxodIK2t8OnlpKw1SjZLvPHkDEv2afxH1HGPPjtUJaT9kRd0sSxeZ4Cuov
/GdK1HSzRiFjDCgIZZf7pHXsDH1m/qlCf3SuDoxbHbbLSjPX5SBwnTNkG+zvpzdyKUcYCxlVEGET
uBpGDl9ivM4xNJSvhrPTBs0r1T6oqrEaDQABYbNbCzPpI8kDUQwU0lLVIkmKGtUbRCcSh3YnqrmW
ZhBFSkINsENHTevJeZkgr+xMTsDc+T6Z3rxxPn0shSrCP844g9A3eLDhXg/X8AuJJZ44ghpUpiTS
XAmRrJogo5/6S9r2FeO6Cn1hgHQ/wRx//je9Lzj9b6z42Ph2m/G7wtpPbyRYao+MzxoO3H9pSR6K
YlcUiOZv52M5TYzaPSjO/zfXi2KE/bvTLPGg5JcOAL9GKpFShxYVV0+MdxPzbvumPRuoSEem/Di9
yZEFKsXoiAep97o66uZw3qOs/qmCNYkLe5Hjd6Kr05qEv9zHurUeeDGmBQl4Z+co7wtjeaL6j5na
rNKkM+E1EWU6rBaHyYRWvMIhA+y9qtqX8wSEfO49aSAWQ7PMKbpTuKfG57AL2/UTfd109uHXoFZw
j+qX/WkzLuzpL+/gzX3gNrKdqIv8noLg0XD0viXquz9uKh1+5aLfmxQwqM9rmeqjep2UKqekOeAz
JG0+Oa3Wz/cyD5b3J347Hye2XvxzcixSzQEX71nKu24E18keXcLhacqUdkhSLR2qTHSEVc1B/xVn
jvtd4Dg8WJCNsymHfywNXQWmHx8Akqqo9l+VehTvXg6XQZQ8r5plWecfpPbABbIBYrZUnvRJ2DKF
OudzF6Ut6v063mDwqptMhkcYBQgWoBUM1HNz/51O66j0hMqCLGkGERBT1nrvqcuR3SZErRwK8jUe
BvcrXqSoBa+KtAdqAKlPi88xbd+RjYgFRz+gBIOqwZRsjNeqQ8hzULqC34l823SwCrt3AOzZfMo7
iaZcXd20gyOh2Od+YZqV3hhr6QwUlpIO51YVtxlVflFypUIQg1Tn/X7iq3rCP5lJzFYd2Cv1ctey
yJ6slvz0VYSYXeJphoJQfJ9JjNHhjYPftqpfbcz4lN3pfoALbfYf94uNTA0KDhXyNOm+X9y+Btnb
gazLvWWUgV3sFVSk7eUTmsDI7WzknREyks5rSkmbSxAGKpSUhsZts95HABBa0LJ5djO329x/HE7Q
pUBEMJlIGns+4VcRgUom9iK8JWqjkMzA0AbEd2i5+kG4H8k/2DZkBFF28B4fWd9n3rwynMpB+czZ
AX6J1Lku0ePByGUK3tTLQ9WH4TkDIHMEUPS/AGz7uV7nJ6zCrNI33Icm1WUnxjsm3JVYX/4LkWow
wyD17epoZZEr2b7tEAxHtowSTVngy8mUM4xRy1eB1lCfoRJQLMp2fpuaCRxyFJcXCZyKrMOoPZcb
fo3FE74HO/WbdjzniCL79iaoZhYnVdCpo81ro5FjR0uWSJz+5Y0gpsWaQozDFM3BxFFz5Z/S+Dyb
SchalaBjdB/v34o6ffqSt53vPAc1jS8LuTQ5RcvYtJUd1uhIcz+T+1FBYvYnX2a4qOqX4ppWWScM
Zu+J7cV88/ipSHR1KLxPLy2oKmmMGvx4/wWqozItL7PLxTtu6vHdDwFhY5vO82VXV1saC719smsB
W399Tplz/DbOn+bSaFNj+tV8ws/Gg5wsLB+RLfV3Web1TaS9L4nHMguI3SKiCmlXTSYNgqGFMVEE
d0GjeQYHyHF89EMteDYTdnxrlv/eWA3lQ8F/wBv97A4ibT1rdDGbKa/Sfo5V3+8cGulBnbrwaKN5
4y9awc3pjc61m2uOnfxhgKWJCHORx6Ohlq+jmeDV+c3w4KyENNoYGBDIuWkAjKRKSPJ2ujjUBHk/
vxU/i36cTo3MtnxmTrQ9JN9CeCQE1lkqIYzLZFAiXERQ+YLBaFGhhTUhGM/edhwipmvszdV+fDQe
qMSwO10jqFvXoeW49dR+IWzXgaQ23s3iAHF87sTcdTR11vyey0VDU8O0f5YgJEZwPnMJ4oGwMqLo
KezV4Hk/k/22Rl7v+yknKaCjLFSF5ntfuM+uFBYpMYAtwU89ODxJ2LDJm5Fbc8224iKr9a7MlOxc
/BrU2xykSacuR+Hw7qLBEdMZogE+buYbfOUw+Whbn7i/lc9KJ0HheKqilbze7q6EzvI0JoBmpIOj
EEME8VMh45JnfHs33koOQLqEEKqLrkrqtyqjCQ8JRYtrZfwfiVaBePYEjYlorxkN50RnL4tAylgj
sRxtQ32RxUJwkwv1tqsk/ejlzzsZ0b4bNNX2Tdl/0Lr+jBlQN4LMH3XsWnXEiZm3crEi/Qv25cBH
F22a1oZxgjmAfJ5s1tEif79kB1CQrFexSwThgK24+Wl0aPAq1sb6cAZX+oBgsVRrY4jBJH48mBiB
+LeGGZVWW5043QmY4X2mpPz9MxcAke1ijuMrnilBwfp+MzyVCRbD1rT71C8KdjNtPxz0yWjMqq3O
3bPMjH3fkR1e0BSP3FqaA2LOWDXxboYU2AbVuhRQCmJlY9TlvJjFjc+k1oMJnOrUJy6eCj1vCT0H
A6CiKN2EQZWmwdP+y1jl2Vl8SBOcJrB80l2/m1BGrofKzXYkd4OJb1+9grWk+yFU271hMgFQhLPJ
nFRku92qSHGTAcGsgydwM1eZoR9qRTavU3OKORkRKgY9aJamX7/5W/6zoRfvCSQvYKHdVlevq9Yf
mmieJ+zK7KlnEBzwe10qZVteSuyiN9h8TDYEmCCwF7iAGnsWdk4SXn+KpTn0D3fpTB0iYRq1dZR9
nKOUbg9sNwMb4tHogksY7j479kSS0qgykLc/fEyArOoNGfnHNXM3WuDzrAbxfsBsQCu7mOSWCFsk
G/vNzIJtWAv9EzVTy7QS4hnlnU3s2k/ZxkqVBMT4hjZpHghCGUxWM9PME1RRcCLuqNs0vzS/vHEf
A6wZ3IermupaHAPmhzeDQ8X1HfNSIyWE9OYyWS0/kO6Pw1MXk6qKeUdjVRtOR8rIb2nYGnfomO8N
y0+kVw2f2dyEaB5TNFWBEhRZBDvOcrh7xQXA9SjCoZ2kJ33FWUnGTRLNdzD9nLJO1W11qEIeTa/o
/oyo3q5FbgVEJ2/u6879YcVxFj4SVLANAAVfAPyx8K9eKLlF/8fir8TrUxyonCj9TCAHw4fEkosf
30J1t+QS/SeB1zfIuw38Ko0nzkDjE6Oh8aY3z81z1UShsQcXFpqabAI8KNHJD0JCatH2dd8tMkde
KFXlGwQYXSBLTs5tig40uuJBqGlnegE4XLlInRHybC8rBPgoIDMslF7kgDzkh0ASVJLdcRKZsko6
JyinVZw9GWoUjmEn5oy13RofMt+wCrsgfymZqGu8pCOpNiHexWHtR2siB2mLXJ5E5VoAToZQoWVW
65yakRoOW1ZTvAIg209Ku9eYfLNzRQRFZEsAF/J6Y4pPT6BfXNvGPkgnxzdGYq1rgPukQO72n21W
HkR07zy5NRzv5i+iR4ApUUc1rEPBeivWVT2+bV27OJ3f1unBDdtlLPb3/dz/qP0nytuGwStMg9Vl
KDGM1NoNYxpBkUNOx6DQjN26hWQQdA7cp9gbugtVt3OskNBBNAeA/l4/dlRokfSWIJLOK9uMs3Na
0gosUuCZErxHJNe8EJ7rnnSUvD4jXzYSNWazImV1oFlg7DFoxeAuNUKM3AmMNh0RZWZ0cmLZjKoP
ESal526MumAUSfT7LygxcIJ/GUzMeUmeVnzp4rLZqHznvn96/oJZXoxD9DNAaGZW+HrePgcXAyet
E1r/zstKSY80a+wR2ilP99wIHOL6wAeacsvDKUHkc6tUhOJJ+KgQFBG1YjRsjk8CNEg6f3W6eF7E
n88EkgW6qCDLniVDAOmHGNTa8KSHTxMA0VzHLQ89XfxG4uL4lhCOnFLP2g+wX9RocP+HimDZlB1k
LMj4KIlISm3eHoug4zRQIan4j5TZ5DB2INg9DAvjTDa0eC/W0BHnVhs5JrOWMWZzG54tSD+25zlx
Ib7t188aEaNd6ai1YmFa3wSu/UK9PRml0a6rdjIym050ubG+JRU8jq2rkI2tcGLLI+890HidatV7
JOiBtpppwO/nchuspCJiF17C5no+dT6TKD9LGajKfvSCdFS6ncQixf/Oy19PZE5FDZDNaUp6yw6S
s4cXtrCkFQ6BkIgrBhFowY7LYVYV7WuPskSHDivjgvUHAGHd9WR3IOho08dHinHLmtVhEhI/NZ7h
zxk8vepazBF82AYsZEDDDVGwWZN6+IWPOe5QTPOc5AHivHSgEHP2IrKytd1rpkowzfZEJEn5YjvE
B+FOcudj9qNH2pcDuQdslwXvUccF27HsKWCHxCNReZLokNsmyHXnGH9Hk/zrzuj7PIYEvQGgzmRF
j3Yrp0Q8UaDfLNBS6m0updcFULccQuirz3RFHtmdyNNrSg40whPKzhHeG4OqRGKN6kctCVZ48ixZ
0/ZrdCG4+HOhuoTvckcm7QKNRCjRls3RXxa9A2noCzCVmcxeKBsxSHGkG2jClaK6eeSf/uQ2NQaN
pMTwsTDKUslHQ83dt0+oJIUZ1l0xlkx4NVqv5PhwGy0R7HQTRNU25I+/PKQV4Wv6rWuIuqILT2Rc
ogeuar3PNDNG2ONsr1fBNrnMAcYqOyh4fboOuEDf+6ANcOw6c0JHwaQ/i5pnTxiGkheTfFFipQoq
Jvi+1QYcNAbosLilwaWB7FqWZYj9vzyIQ+Gv0u4jZaSoY73wUyI4ThO/MjntzzWOYseZO9lD+3vy
ynbbQKrx2C6mccuzwOwzjrrg4Gr49Dx5GbnNiIkHTGq7C88LNSms1LjdiwF0xRZvm0GiYeMZ4rdM
vXqNYYdlvmihn75u8d9nlkh4DOqKRxP/yaFShtdbDkumVU0OKu6DtpntCLuHfqHMdmDimfz4cKWZ
FMZ1Ml1dnZwmQI+ROBCF2Q1wZYH7aLA0gO9hQ6EAHrK6ZwOCUMUGpJq7mISPXu3SkIG/4TKtGspv
+fO14V8gcdqB1KiHNqRaiMMkPO6I9ABltcHOONEkg0FHulPE4V2ZNNK/g2bdBtbvoxtk2sEwVBEH
9HEXSVbpWURiv19Pv3cYjw8CgEbQYlZvrayxqI8/MeXQgW2wQcW8xSsHoP253Glmydan5WcqYEEs
kEQXE5UpdUES0vfnmj7wM32sAMdWNp4qwXLphxBtVOfQK9KDdfKYtJ77fRy34vIadOlp9D8W4Glp
Q2a/b+33XWiyzKXm9f0qOEDe7/7nE08DvxdwiXHx/5WCi1HL0CFtAn82PeANRVEiuuZpdVhrOC12
46NGTq4skZx1AkedaLfu+hEC+0+lLtQ5qyz5MJHkSipGxggtsSRoHb8H8WXHMedyt7A1AK2be2Zm
LEvSRMIeJyAJXz6mXSdFp8Lbl2vfj1IKCVbNVy+gTBA9LyTcQ1YVU5I6Vq+Wncefv0vRRKj0auEg
/qFAwYV/8Kp6czOO317Vqkn/D2jvOQX3+1cvEdILZz/UmhqBuwPPu/ghWoilrwk0KFwpleNIII3Y
vqY09uGQ6x3qUE7fhHdGKaWF3sp7uf2m5+qkxWMaKE0thqjQ7jMlll1Ms0SLTI/4NPyGVOUPmAhC
tYD4Nfdub0izigoemNdF0GzZepjODTVS8G4GtoG6sYXqOwSspahXisJjL+4ZtDlS5E95oTxDouzA
AODpfPqY7vKYYdXxAloBUe1qq0fuwHFvyq08Rw4u88B4XJYiAvb+9qN6nTa+zop4LAxtgrQ87BSO
BciiTUPAc3WfPTPG114Oje0Bht2vPhZGoJ8TA0Lbsex0ZyRgfTIwbO96d9v5J1TI2WkmEynVyZ2H
qTDhy7flS41c92zYtZzxweSuzEbbDU2/0YlY9rHnlFtjJrgBZzmG0Rzj1LIzzkNb+QEtkdnHBTRl
96V2tn5GRFrDHf++rYxUJHjvGaAbEm73w4YDvm0XHdE/XeImye2nO6T003yDv+8qzmMFo937K17U
PrVWa2EJ6m+9sWvVyy3eGmdyc8/6Z+vReYNI09CnuF4gL20QevznfiJOg53CaXnm/PUjAX4HLTXn
8AgcAhAABJDyC8k/Gt3r4TQsCcWx9u6FpIQpqa3wi4NxSG6uByUzstl3poSBnlHaWi85Y1SFKX2W
qBsMa5hCmoGYMQtfG0+UcTabYqPYwbMoSg8kvT5tscSYCFFWN3RfVmcqLIcNPj0hK6Vl4uL4HI8l
L89cCy3msxjIXstrT75B4XsUKtIuPWoD8/kZFRUMkFP5dhDCpIre5lJQ/bTctV4IKWeNxAvOtfZp
2jJLtPvnqpGDGk2wrvJ8oD1HHJka5pm8ev2dQ6j0eYM9qApLXD4qlKgaOUZekNynRrta0/H6N1Ft
nM3hhZsY9ywQH+TlyTqL0wLQA4XPpGvUasP1moDLgkh/bI3OTdifVhuqAV0MNpRIAh4AadO6FiuS
fYG8XZvQcNcfhxdzKD5YQTgT/C0PHp7Itfu8qlRE6+cC82kjBPHs3KNDraDjFJzHHvvimT9VtXG/
Crydd4u0B3F0ZvusjLxveejtfGeuMwGD4J4GI9zaEzAy/OkN6BxKpHquTDlycx0SZGXuHItRj8Uq
wC9yqOrUnOv/kJdNE6ONB9bxl56/k6DliiStghFkV4b0IkV5M6frA5h1ycxCCE6FbsNe3hSNuczG
HeAej50Pm5jUXtcs2ZSK1sFIx0hJLQTCUWsqkvnLa8apT+pr0hIs6m6Vh6QZWJ6nJzcvJpyihw8I
j2rwhoQLAC2HysPaqXuv5QPqliskhobVuqYA5D3udxc/eyOLQizhfG3yPuxTLMvS4UENwRqgb7Ld
LMW5uYoZ9PErUQg1y1b79S0BGxXer1EITfEH9CM4py5e3HRC9/pD5wilizTdNGxFPeyB5M3rjoO6
uEZ4RjpIifmUoxGIpyDvrav3onJerLiRs5+QkvSkYwdnFY53UPs/SUiaBQhIHuKMeArn/Q10Rgae
u5Mm0FZCVriig0zgZPq+hnwF2CFfYBmJR52+HNFOQWHEWL0Brok+TKO1CyYrCG/FOU8UNCtGbKEI
VKfDi56N8mEBDlaUJOJ6uGzsX5llVF/zYtnaJIAJj49vnPit9piQeDAJd3yP9v5q5p9RYUYSmOko
Vu/5EhdOcLwPRgBE+SIog7dH5y5AT3yv8HgKs5RWy1dS+m4HCAcCFzCO5USUxrCkK6nVTYqUE1X6
RBLE7E8Qm88GRGHq1HoAGQJQOxgV+CVSquMChLNsIIpQPgw1JuSuxsPZjUqqGt5o44hFeTIV5sJv
IVtsYDoYERJKEI3kg69Po0SRr3dqhZAq4bOe0gYHIX7ISUzCUlzg6gZlGuFouCTUypvHfFTzx7L7
1bgp0vnoEr+sS9/xTsw7RmNcroQQZaf3AAH+rEV9H3w6hR81vo2iGJynGP+IvUn+zRPtzRyCzBo9
GsVrGo3J25tNkPgF8DLdXemCWCVkNKjSTuL9NEYuk4ScHACQbDPivG01sQM4xgkMvDsip4+HSZ+d
7IsqmqRbvJ/HrZk+LKWqQm+N5jsn37O70y3sEdvKbQr6y6GA8wFSdUKA7f1FpzllUAjitiSlbkfz
da7ic6GXD3RMS+K1RmSDEQOtEFZSgRGTI3/SwgI5F2kGaVKWf3Z4B5VNFiKHuvHlsTC8bmRKb74H
9RnzXhseaX7JYgYRoSeeLAr8edlif9FQQwn+LkqfEcbaQi6OoYN8BpZ82X3m+bdNyxNahNX59pUc
LebJtie0fVqE+Voaq1EXe/kii7tDvw5zVVIHPmyoSjHvsynigfDDvTkOARUlU0UbWg8hRuHYQ+D/
9AADD6LEQoLfOsSNqDWnzZLn+NhPL0By8eO2DmTO+l6Lr+PV1emGshuvQPJuktkLdBK9qKwKVilw
jrew49upMg5iqdA1A4+5SBNqzrmZTvixvUvp6fAhtNVYhC3ilrSDTgSoI6ejBJBtazJrOGr0swDs
aMUHMPR4FXTpnsM3mtQQNJmzxtbvNSni42lWkzLQP/Jjcyz07r5I9Lj3eZGt3xwbo0eILRXe5gMI
5zklf1h3vsN1svnBpxE8r6qPJUyZiknJC/TysBFajeuzKEGrPrcruQ8Yydnke3qIYQvOjG+D6/vf
jMphoOOQr9dESGQnKP94765Ogh08GSIV7EFvAYXiGPtJ03Yte428EJbxyte1u+LWwfUW4CcJywRV
m0zlVVVYnNTTbMNGyVatFR4D1NgcRkGD3tUpTK1TsWHwUGtym7tECeH11EUMZw2CBYHbCG/W8RP+
FQ76T31xxNs73rKoqKahsDIhnpJB3eqaDRATcAPygEKgVKGBNUOQZtAyOiKDEGmgX3KCwhfbxAjW
nR6FMJjW4ebKyryBS2hqujsxy9pw4pMk1wurWBZfvFY9iO/2w5yB3Qlz/zvolDNy7O61bd9N3PvY
Zt24rR2907+A9EZrbLD0XcU5g6XXu/4tQrKx2EmgHlPRuXHfqzn3if++sewgcoFKYGMYCjSvjg9o
V2RFBpcv+FLkDBEFW+N6Tk1Al90xtRbYt+lk1HY9elAhYCMHCAVSPYPY1xokr2ehDvXqol9CxcMC
0gyXIr5pT9bfNNVJykNLX9K786vG9HN6rvjNj17XVLMehzj/NQtMrOp3/d0i7ljU7R3KW5UTMRpa
VUJ7rFI9oPYe+rBYSywLLXFfDYVH/P8AqcAIHfAJr8ewqvUwn4WE3Tf7JvdU6gDGU2JEBryz1nhm
DCL+6nzNHiO/Us7VKJ4Yc+GKtUlvi27J1ux5CheJjTBwfEywEFXYwvBych4Hy7UrEbkjvBZvUqq9
OcRaOFDrkcTQc1DyGaWd/JaFiAhjcRCBGyfNgXVeNlITzQ4xOkk8qQA2p4tJYHEASLK8uneVavv9
5CfzGUcxl0E5bpJDFFOzW+Tjvot/Z5tWI9yI4nBJQSEMry9m6+HSZrix4ipadCs2/O5WJOs1RB25
eIfItTVFG6A2G8J7wvws3bq/yww6RzZREYfWasoZFgzvrm1NH5MrrM8odvnVuEi0Fbh8uPRQTuRd
h9YVC6XFQs9Ej82QBw5l3ZmKWlQBpj4f3q8BaKIlvUJGABnVR8XigR7RwbXY88HLGJN1bG4K1xul
n//J85HR90hDiURkpw/3nCMnALWClTRFRCWueQodCbq8dGvFgqYcaahW8h1e6EkpzRhUDD9gyDH6
Tat/V+e20R9hYmie7RNoOBCSBhEAs3QNdV8DuR/F/O95FYIMp9SzozQehP7c5nAWPgwOe/Mezovl
m5loNsxRbnJRy565Rqgl4IxT6JJ7qS6OTiguDgKidzHuw30XasyKbNTbJoE2qy4QpLY0usFVtJuF
e8R5bdJHHgDZymDTPS/2ZOxYoP9Lr0Jp3V2QFFYQfjNXgce0R3AP/o04QnEY2C0ipvPvcCS8Ja88
zmQQ/joQQ7JPKlqDwRuyzi52+P/2KM2uY3kfrM74/bMoJeiSt54u9t++V+8e421OhhF1KpaiCrWi
eH5yZJe/qnOgcUKwKSFhcUsQbrCtyddtKhROtG4DiC66xHDt2tcn0cY99cIKv+GSsYFZt85UWL2P
/TjX+4PJHsh/aLOugan+NYR13lMkYK2x+k2OtRnA9Aok5GKvU8dSUVh64by3q4PEw0Ee/tT7hLMj
v1XQU4AtyuLpfQswV2LJ0d1d3QAzm/VNNkQWBmlb5hdHkzY+Us6ShJBmQ367GXS8nU4kF4cQ5mqU
D+bp1fSgSj5ngrH6JJXbnmNxAcGyOgG7U/5MMAWCarSHD6NFwwyA6bgGKclNsaX6U3E2SdoTV5Va
ou99ueimqMlwYbHXwhVlokarZPOh8lqY89z+KteSnIMziTVHpavd6UaS9TeM5dXQFjtClVgfUYRF
yhOye7ASgg7M3MBCOhq8gvx7V5iKP/giMca+jMYQ+aA7xiyRboP0OTd5icyXJpkRV1jpC5065dBA
9We/xpZWk8dS1bymFWFO6r3BfHiy7W+cSG4Ncg1Qpu6wLUDH1MVwCQq8h5709LrDjfZ/lLDBuc9W
GoSLCa5WtHrCrC+WZ6JnaVIiu5cZ3c+GPqBJJumqPc+w0c355klvyRSzq057smM/N1t+bkBVpMoz
0r2EcufQ7T1VkzbC1Yb1ZzHpz6ank4FaMhEkpYDwNeZjrHDBNGqaqonUMi1fhaIdnNJnvAGJW4dc
PCXv1mllVPVOLLGXtgyN0FZX+gAZTZJIfIVODrXlykReNtNFw03DcRV8wtYN0KZ1Ev+5S8R3CA0A
2suqZ/M5hzcvpX/zkTnSBFHnnCfkcE6BYVc1bigIFJNmcwisj379jcb5sVRMUXulKEOTl7MdT8MZ
CGdAAAGQQkyJl0/e0V7/sgQpGXjnD8eNpJo7m6S+yu42x09414FKtr0Yz2bv8mpacx+gDkMAe3A2
un73c/iosaOhq6ffWeu9Qh1sb8maI79GPF6nFa2aFLTRPkRxk3HalQNMbvurtgf0HR9P2QtD6/33
px2yDwu3eNUL2BHvfPoAPYdbzZFPLxz3X5eK9lwBBEjqTLUzlwSAf8PHT2orpSw+SRgfZTqwUy8/
VRLU6b2x217n0DlmuI//stN25C+UATqsnFzT/q19dmgMMEf+/CKeCXFXgtIPUDh1p4uM2nmdhLVE
CsAlTZ307bOPogRTw/ypWHwnhVsGlET9bTnS3FDsAnXfrIKwgCIlLCHqmBvQZvpzRnMSs+lY+tsn
BRy9EAI6NLxcvdlKYbErgv3qNY6wmajHzfqNmPxD5sr0pRpGTDN1QB7Z665GEmj+BbTNp7iTkpQ3
za/U4UtwLbOtzb50YNxxLyzslRh0x+Js8MFKiPe2XPMHYEhjlE+YohOIWfC8fLQ9puRW9+gVO2LR
BLZcjYguPSxu+y6ltNneZ09t6bY167DAfH9D5rzTGakLVSoGGs5BFUO9iRn1X001SNWkpF/mOdu0
vO3IKEF+TmABi2FzKGiYp7otCRBm70jsjE+L2Z9qq3oZs39kvIsOJ+t1TBJzkzHdX/J2n+oXEJlS
kN6HkxNuEInxG9nA2vC+s6rHo+89anWnu+zOKh1/uxxjW/G1eNXL6OyYnEOm8qrRnODRsQEpdrow
5HoiLye5S+g47nxaZQHGXf1eDbigyzgTPyi1lLxEBBh78P94Rl9rJ9GH4/7JJg9ZLNRzZLLPJ1iO
DNhQ6qvXPu/Gs/3gR6aibx/bksKPBCb6rPvVzQv+dUKxcVn3tC3Mx5j3hnpj2YxBOHY6Si20Khfh
NU8124o65qQWke7T7E/Lkpw0rgR8Gw/4i5Kfxi82EmUZqCHwLaBWvwyAMzF2LKMH0Cvq3wCM1QPE
Ya0wgtUoV1bKuFalpD/V79ccFbOfSsJRD1KjuNJmOuxUllqhccT6lxrbZhHijVCYmQySezgXbVtX
mc/3LhAXgXrCUq59hC+2FX1cA70CPoZDfNSVyZ7nTDeVf3NwNyQYsuQyg38vgI3+/h0ezzuufJjc
kIMcA+0WWdS4OlFhRhW62HqJ9cZvowZminCw3MRan631w2nB4kp5K6mwclREkAcOZQT3KhOrEMju
h+wzt4ZYPv0fzsaKvFcayDszlI7b08ccdY3f/N25x4NV6tUlm1EROw+tzqqQ2B3CTEEvHlf1YNiQ
t0cbsKqTXZWu4hkObIBhIuhLJYWsnTH9d1aflkOeXgaPNCot1xO3MtTjPTwzL+VcqdTKi/VAd8XP
Vd9AoQxZ7/uTTowdOiFSzia4NTINFetMiF43kj3dbr4EOZ1aTG3ti6OQB3pnfKaj9xejlIx9XX+k
3J8zP9sI7CG/pZYMDr4ui8WqAhUMQjo67+SQ9b2hjizKZQWz683Rddf4WK4zmuXUn22T9jQxvrar
KX+HDpx6J8uOjCiionzECAoSMujOJxQdXc//m4nx/WgqeJsuxMaofxxqNTHqZd9k+q881X/WTur0
v7EhpDyQAGCZ78oIas2Z39xGjIMPl6Jumz26OSPh0g0vPmGb9hNItQSbO3jJI4mZfmi6/6BChhbE
NzBu4BHFuuy+3tGoW9cZXO35HE0CKLXUz45mpYJ8VP0XPS7ShXesGidIfF2FBbIAUu8+aMC1QAo3
wNMFZ2HL0ro6rzpOltNxSB9pA1I2PzyBLKu+VZwr5DlkT92jA1l3hUd8oTy8JnnqENJ5uLQh3Au/
Qi7r01+TY1EtxMlvw7+b0euTX8u8feNLf72gL7++URvEvNzplagh7bGLSSc4NoDkQW3NQsWsNRu9
55AB3zYyJyE97arF9Mygo12YYVTdVl4c+OdizK2EtX0OwZURyCJEv4+yjRMnzHPiPvfb24ier2Cm
g+2zajtFWYNeKr+t57+LiNQYSLJLKRX8N4mI6vnERunqUgpBVhDecvmW5irnrC1bwbyjbCr2u9oT
k5xElzL7rLKFyqam9SzZymyjobSIcToHnakpig4311A/SOPXzto2fvpx0FhXms3BYZU+dPN4THF0
WIaHUb29OxjvkXCTRLEH2GFmjP0OpA4tVfhazwYM570soTnPpQjhQItK8uPf/t+SsW9CleI/w/os
bqbpJGMfOl0oAo/T/s3SD0B1fMCcwoZJDLTBjF3OK2TG6nlXCesON/uxhNKwC9bOvc5Z/PlJfqFl
E0raPnwbCkh3/n6A9DyU3qwxvhmTOGVNKdiwgiKL/vZc+yCCi/sIqBtWKW8wvPAfOccRo5Wz298f
tvtE0Yi6CeBxKJLqynf/QHx5lMw0MsU/b9XCyT7XxW993vxfXJF9rLtcm3BfbAc8SplbGhZCzrrS
PzxVQZVaU3aI3IwobCSgZ/6lNi4Wg3DxHnlSWgwvLV8L29Ln9czjE6PLZlKIc6gQ2cUbgTXVhwXC
kEW1YDl0+z0ueQWbXevx4O7jOI7sQuz9ej138bWK4fVO60dEnPcCK77ym9ua5DJWiBBxMLAgRwGC
zpX/0DFRXDXeCAuBLI1z+OAc2t4+8XjhfxWzsrrau+g/HJb+wQU/BNaJJfDS+FMs+6FDMYlZyn58
qHaFm5HIy/XgpAT30vUBPXeEDEE/3jzPgLzLx4tXPb6mc0pk/0g4a5nDokhVJkPOp9n/FPKow1P/
aizeXRJUm7OhOuvyZCHHvsO8SlFgMNJAaollzUaKSnSHBI5Vi6r1mfwcTCgtvbE/GAAHfk361JYc
njWzB30Rf4cRNyDKFH+lI7cDZ5z9MQAqAHaoSu71GajcGlZoxYjiHosS5GGBCZw451WONplMyE22
HtnSLVyMKkwwrKpR5qtDLpvnxU5tO1xejyZ5SYNcualTIUmZB6xbyU8/3Xy2Ep8QOlcUBEyQw14j
BtBnxRO9uW7MheUDq5+H3Nnxo7grwUCWp+NalycGV/p+cb9+PJUpBvOfLq/VT3eCboIkNNBMKm7/
eH4Kwy8wWiLLvq3S7M+V1L6NQzm0pWkFLQrXZm1B673lc5VjI6hV9kPip2yuhbHl9L+Ezmy8jQxI
IzVJkLYAMhQ1GjYO0ZTpQgN/ZSU70U40eOP33J2h+Gix95CQzcwdEUbgqu3WgkFIcDNg/Tz6OVGf
lLRG8CZpkccU2OFxYtAvIq5M8uOC6gB6uColNjsBIYfdc7ys1oJTj0lpi79VzO8wCVScys2mJpg2
7scJj8eYEQFznjcQexZOOMljBuk4FwIIaarkGX3eLctqzx4nRiwifrClu3KHZGShMcYIiGUfGYJ3
UBMqyY+vet8RuolulxMO8rANgqCuZFsInyaUulD6ATRxXfVQlBgdW8slFU4yKQDk2LsVUxqAE/iV
UoTPPAiy13l0f+r+0nFk71mqmjqg3P8kbxnGJRl7CC/GzHuBlAKPlvsI6Vkd7agnumh1lOwCJILn
bwUupstTmrtz8D21768JUtg3Rr2QfK9ot/jiFdr5Piq4f4IWgHo4hyWJtzrALuH/iH6V3Gs8hTy0
1+GDlmD0T0b947NARvlFKtUr0cuKLIhZplGeZYeqBznPrFDeUr4Ev7IuWiMAkT/wIslMy6FBrgVO
+qCvqtJjr5zcUYxHj64Nv4BKikylY7Zrsp0Z08X6Wb5L9MY1ARiAK3EjkDBklefKSuDV1t4qZJby
hpeEM6TQZvlm2VYGaT91hy/5ug5nDO9w6JlI3tW3MGsnfTikCcVrNKVV9mN5qEDeV0VMoiewLUzK
mKnItD6SH9Kvu2dOkRcx/CJjOl8pbOzTmr2xMaElIZjdUznmJiR0RtMt3montjtWSZXCyLcDwq9P
lDtE8dlunOdOURuuz9MWJGqk/m55CGBE8SWnkeyd2SqbV0kJW9ycaeI1XyqJ7IU0JKLd/EKLohsW
mA1Dx3o5VEO/AJNq6NhjUC1WwCLVEgr8fuVTTK+GzyNi7oCSLnzrdoTrBhw1EGgCKCDJjZe19iS4
FIeyF+AxDpA0OcK6lnxgRc2BELo9qVX3aMyPcIXH1nbSZ5/SYVUAhki7i9MSHm99Wm8Bevxss413
sdGVI/Ft8afpYbG+irOF69bO8UGViZyyundfRYDrvDY6labyaEuRnWyHHlUf+nL8lK7oGoH5I67U
TjxC1mVEo6q5PaDso+3CjNA0khLua0RC1WvC/mxbC4tinFjzhPh0UPrymy9hsteGOgMcF4aMPKns
AG5+QtVtMbrUt3pYb+3Jt2ZuiU740T5zPgb4Vftvm33aw5m6ewqJylIEw5YLIvn/SBrkLkmJLtgc
Yt6GZTpruugv0haBxm/QrUUt0th9LH2AGOWsS6FCtL8APRS1RdNcZYvdarbSND7EyuVPSHai18pF
4sn61f3NwjIhgw2+yz3I1yC7I5R4MH37vuhaU+gmxSl8XRzUwKj7HeCm2ghUNt6T8bDlHXpC0Fah
c9N827XFBR8UE2Hlc6HFUWlf2Igsp/1NNRcblaiFBzpNcUmBOQOdyfTJjAWqrVP2quptmZFT4z47
dDhRVM2rjjWfhrzPniPAz9jUBrhEvqjVrqrpnv7pWmIl+m7e/AsxKqW+RoKQ2g812aNxx3qs/dzy
A/TNaV6mj+qaiKEaZ5TP5RNiJAJM3fnp30NNHPvhbtV6NPi9yXAlsGUIDrb+Bb2DLCxXPqVUInUU
ILVURw7GADZh8m2o+vlJzYTK4gFUPW7QFXCuBR024TXvZEB+JGm/ROVv7s0Gqf8Nsz3CLSC8HCHZ
n8Ple2qKb7mkFmHVIs7p+z1i80zoDvYZUdY7NR26+fGU4OtZlfSom1nmhrirBEJ8yNjJ73KdqlqD
3rFn5lFRS3GWtGsvkfYpdHeqQyi0DHzieVsAcbJS55Y+eLKJaAGDSJUYJdsrJ2P4BaG6JWN1q67H
oMzJDKmDw8Z/bBVK6S23N/SByWaaHUpXygyHfD8eIQCZUC9wmyoOKwc0rtnrDf5RMoPevmZhobVO
01yoQanH/JuQ5uYiAzWHsAMxpN4/4KZR0YFZqJwZYaABxl+2u957R3dN6nx/Gp4D39Jh14nBERob
Xx56MS3UD+YguIqZHxONe03Y26uvFuhrWtPeWgkJMOlUB60SB1j4UABKWqMJg2KXMRWCQHpHYoyl
8cYMDRmBsXjEyAV6TCJ82ub5IObGVsBqKN+6TEv/hDqwCQWJcGEHBLnvwLYgPLquWvSh36a4HONM
Ju8TZ6xOjnm3GjvmhkljdrG6p3Q6dCLM33iuCTwn0KtD2miLUZ0wPokhDheeuHno7SftoUljDSdr
Mr+qE4h/wkkal1Hlcdh+CaGROMclr2i+AkzBkWwZBFN61pdH+N108/rZvW5W5LNdbhZDSAj0NhTg
EEfD+k2ve/jPXMpXRhX7cG2rhn0AGC6FNJiXV0Nr2cZql3zEOPgaXL8DnVtmmhwmxAG+2XnajKbl
feN7qNfQCXhdNVB42ByGVVHF3JwWpDNRjX3lY5oWbieSUDAsY//0WEi8Oh30x0tdw6EolX2VpM2Y
kvWy7hLdaRqRdyreGO+h7bnb5TkZf/GPH9NF/m/fCJLyB+UbI919Yqg8cSxoURuq9L40B8Tg6tCN
bXe+cKw3rjFWZp09nxDinNwFRSOyYtzl53hsvwsnRpPNvm278FW7wwsH74fH+842JHWizMRHeqBp
CBUqAdww5/E+DqRxve50Vn2TuoGRbDJ4FIGw6cMki6kBlio8ccBAMn6c0DR9pXiNjEguB0zPaWTF
2ritpXPB4Z8eFZTCC+cYexRt03ItVxIbRdLU2NYQh5kRHyZFkpKOtNczHDTCBdUeWNFS/R7PcAV9
KB0JjEqoq35IextqOXFcau68TDf607Aj2CvI6oArAbYLSbM/WpsDg3wTMWojHN9frM0fAd98MvEX
1r6c8wyrO9S6qsvHnnWd59eNzSqXiayUA2EQzaK8dIe1L4twMp17AdRaxxL1RMFm57xNirn3JT0Y
EwxygOU5kMGWoidOHhyC63/YSbyIfnEwpV1bY1eFbbV2Cw1r8tU8R8DO/NS4/GzwGoFxLwH7yBkX
fJrMK7i6XBC/9O+vtC3VSVZPKyFdyKtlLl7prC3YQu5Or4vlYIg5C4+F8opIuWlubvDf9kyafwYj
x+p+e6DC8t137GKg0a2rpH6NadrVYlUe75VZVZasO2Iu7Ug6qRJU/8pyJSrWmB1lNrpL4nge4K+o
q9A7ozUM4POdB/PjYT43+oP4eujxFl6yzX45k69Rw9c9msGyBB8HWF30VuD6IRuSKYY/g0GR7HH5
VoDp7Tq9+eLUIuySer6gsVHwEw3QIyORoFyc5pYTeO7wTRk8tSO4vInRyjVPE63WqI/Kpj3LTDdA
rFsxdt1gFS4Ct0/Pox36ttyDK+ItbRpkqq+IiIw+sBaMC8lNWHvoj4YwkoxJVzmRgnfqAPxuBtsx
QMEuSCXo8R7ZQS1qwald45Sh4pgEPcYDF3p5SuEQOAvL33Oj6yA5/+ijs4IQazOW5XMEc189BI/2
0fvujdpg0B4wz/u5t5Hblbqpyiqz3+yza/0AFib5gmGDaE00ckzwdeyMMyEyJDAJcBZqT7Pk13bj
GMov98AiRrQtumyRK9SgeFbA/EybBlSm//sZ6tzcZQ+c50v3scqSGjaqW0EnvKn1iz11C2vs4CoU
9X8XXThK7Q16xbRVrPubDRT8sMjtqCZHRQ+wHwxiW53GdFU9MBtyPkYAzg3M4BczUppcU/wTN2JX
iLN8We40yKQ+W6AYUN36zLKP24/xdH/Lwy/kL2YDKAriOfEDQxifZNb98EN4zjock4ngadzn+Gbm
wernXuYFO+3zIebDH+DoglBBOd3WUEQyEgSIyNXi/OZWIvxM4qpWOMO3CUz4P22Eg5n9xfTC6dXx
ObAlZwSJEkFVpinUieAbdEJ+Kd3kDWCnN6/ggm2J/XKe7fpb+IRgcWoK6lW8GITrVuGhsHxXC96p
/5PPy6SELLtOPzsz0WMVOT5PCNkC8vN0h8omRwXkwBHvBSF9LCPnd+EnAlHPSTOlYAfaIG1miQxZ
sKy0gr7Y5vc2f4WWDyrNYZlhw0hH3dNRJE2OBJVSbiVqc39FUuBYsBUUCOtPWD+Dvq5HTAnQXn1f
3q16XnUNDrifW0PYsauUcmj6eU1fVFItgGHQHdxPN3osxEY9HwFZzn8tSTdM5FkRO1doS2rpa6hC
SpA3PcA2MEow0nx7TBfOQGyk/HK+OAlQLP4REqnlVUCJjB25pWaYxsiMBYepM+LDfcJF9UlOxYoM
WxStjgcaNqmvGlTmqoiH8ovp5ZkMbbz8lWDf1zM1iXePd7vsVDl4OoZBg+BSiyPjZqWayTgD0TDD
UHwzr09DeodXsGTS6sArEbliDbn2q+cCu8I019rd/O7chSc5l+unSdq1rgX+Tixqz/Oc16Eupp6+
IcknYkxlk2ES2CVLzaKnPeJ3AciudSYAX0YfDOyOqUMBMZZT7Kg/n7DyXuiNt+jXcHLpKnzO91N6
/X2knnTO/e35+eN3gPxLRIaedPuEzWC/p6ilVqrG7o8+uBiGYjbXns22p4SzwA1B0984TraPVhwq
zNxiM2cP8+R/u1u14XgrnwhjdsY67LaaGSQ4QVJ/nJaV+qplSfuQcz208FM2p/uxHaHew9S5+P65
kO/Ql1ktsJHkJTz8lQZQ/PXz3BQqJG+FRfBdoFCrYOmzZj4fJu93ZrbSCaFj+UMDb4Or4UMPd5aV
/XmaWcOOeQsJJ3CDF8TJtIXj8CHFMEUFcKdmQQ4L8u4t5VWm5I+j6kE2C/UXXCsMaz9mWibUM6hv
cs42RpmM9KumgW9EfOQz1Na4P4GJOo2DcgnOZrm5xhOtFpF/lus5SQlyP4kx/58zxxv3A9gEXCZi
MfsnYYGQneKTOqSpo9keHYz8eKEGR/MUmPrikphZwV+myTex9IwLDiLZt+lTnIP0ArzTw5IJ8nfS
IVuyJZ+vGrz6BPUpApeQj3yElGBUOtigWSmon5nF0m9f5sORvgsc3NSWPzli80re5fM2eIJRz0aZ
h6Sz93pUl3p85seszR0YHmat88Q54BYtCcKY1gmtHFM3WKiQW9Nv14H4MxsQPtJjkbtyaW1Tohzj
khdgKPVcWA/xDJU0yl+L+l5DAODkhmwnMrtFgK/3vMIxWQgl49ZMuLwoN28c2jAHGWD5xVoZbxPf
fDSzDFaJd51+yjQ/YbK9zVxBVnbR825tcgiPvk6s1JgpRxtRsOyB3QEk2zjNmme0GvU+Ltuv+nJv
XraPf0HXcuOmNooaL0ZF4G5675qcM9nGhgqX6+rvcQ7bbujkuDWNrJXlS1H6XPMv6glR1a6eFiRr
qw7Nh54fYkSRIkTjt76W1uRXsnkdPBrE7pdo4GAtmBx8jsHHpkZJZki20Vv5gcXuRaUBc5jLw3HS
11VvMqk39GIS2qIpsNuJaIce6ozG82WZOXmh2hyWMznIfl1cWI7prq5/z0FaCCsRNuEbUaXBYW3K
NtvNee/DPHCuC7ANWyEzVKmMetO6MAc++wuO7oF0F7b6wzgwuoZhlr0CBIR0mI0enaKdeg9Q0eFx
euadyPyeSzzDq3arXDHi7UPoMUlVhHDnKBRDf9p2wVVgihAAffhBLeDmqt5MAS/nHyKpzaahsGR8
5bp4boiMicAEZzhkWiFRlsM44rvQvtM0A11+YK9qPSqavtJzDNesXouHzWM+js9LNOUEDnYBpIvr
RuUQoOnfQwxH+PP/dYSOyqAxZ83NiuRH6BmgSc9DAtcyzq3G2RLOHsYE27eBb8pFwGO8fHJpyjXU
CrhEojzgWQiQc7JikiEVdtUgzed8xJ1xtUubSd0SCwaFzvwTFJqEvJS+3kn/o3SmAs9OgjwedyGu
x9/OiEzUPddKxOkNfsytRihJjk/O/x1siNt1I74p4m5eI+JfmkgSavvyebPFVIZ88ZLcVgzqTE9G
XdFJdhRc/84vK6lIRhO+uCVG2nbqrtCf3H8j+mGr92fCzxbgmZ9K2qd07eCXR1Pe9xNM23PfXRMP
DbC0KqPd2D5iR7B9n0e5QRwwa1qozDkjgu9q1UIWkWDp21R65lVb1hpN7NgvWpHOom8i+jKHC3uq
HiSCkdv7dRKzGDqbqy2Ye2wzVLPTn4lGNqPfvgi/+4zMhJ3v+rqpcsrx3S9/EwBiR82PMkPGN5eI
RTEfIqCHHIOmf8INzpakc+yzqTwJ3+TUwGk5zGy/7n1dmSn+SZrdt/x3NpgnH8WudQC8Q3MCr/wN
a0KjhS/FuCFXhffGKxuuwxDS+Jx1TDIrPCmPD44InRjcI4Oa0iqiuPgwW5tr78oGL4Hu7GW7reX9
vSX7yMBvTDfWbZKuIRspSb+/OW5mWmuIRRj+qY05t+fzt03MIPjSWu1MeIm5dRhaiYkN/sy74yvA
7l07zdr516VXmqz2yDSFSLwUVOGe7nPT68MCkcwad0GY63ZDgots5DOe9zt9kdvy1Q5ObnS4UVra
uRwjP18y431fwKx5PNnMQqvHgHn0m/ky5lLYvBXCrR0zYp53OeftKhq2pl/7dniPyCydXP0eWe0i
iDWEXhpOV7gJUyfxNIAiDLGxzeFbzh4hOD7qZWT6gkGK1eOV/mJIOVsudzeWa1+HWUldjUrDF1ti
uq7IWQ4TIcMWcrE0uWc1q+rHE+rxgOH9j3kuG4hRuyEf06MvZtAzz8ciVRnAIAidlY/nqmgkeCkG
aLjQ55Be4lpJd1Xiuu9vLbnwBARi+M+3+VfVJlLLhxXy9PJmyG+ooBU6LegGK3Q31c+HBlkPZO/H
rog2iLUexTb09fjgIXhV5Sdx5C9Fje49GyRh+ZbyX6VL6eejL/g9i5061zXnneqvQl0kaDWbruhj
XiC6bghTdjHR8PVjA5qQr4Woig2e3VKcsRAS18Mz2CHNir2wR+grA316UXr1WARunaijSrQHFE/Q
HjEv9Z6Wrv2DDOk/3hHY+SR29JDnJi07lI9V2gvTTHrcpelIcTvNWu7BtPXHZ3C8IyJhF+QHz3aP
1U7ys0XK5IUOXDU08Rku/MH7OCWfq0bUrHxjq4cyfiGoH0PYCL3hob8LKfxH3cxHB1HnqD8gplwy
nxJHA0a9wYzEiAAakHYsEYJ2WLvGvowiYSbWGJ7JuuXwBsomcEz2O9IeOnYi2GhA8cuKkJ6QOlnf
usNDBM32Gc99rPnPg+Nb0A5VDV2sZb6ycAN6pFV6VPsGqNm32E86Uoi9sf+s2sgRgb40l2nx5m9h
PVt5xmqr+I6YfGUPdD0FiJiEGLvccbRkiPGl2vaK0HpQ2sR4eN0X9iiI1/r6L9gyl97M92wxivTl
6QAE5Xpmo6qoNgxq5BPFFg0AFZ1crmBaTJeTpIC6Dj33HYvMHtkzueI9PC8I8uhhOKUdZLvaFSNc
ObgJ5fDiibWoxErLiFIWVA7jht/3hVhGDuSR1s4RuTmgCLdBTg8oWgP0tKamK4zokDhlueILxD29
aVjOxhWTjvqIxSLzjVm37Owr0yGbYYWvxS1JlFDt8q5b1pVmWCSL1PjUzz5+kn6b8li0mwaM2kkF
QhXOEMR9N610REmMvvRm8wbTlXxz2rRnKecjkQO34csXggvLOILLSzMoy9sSxv30oWFidqHP3MX7
b7UwOAops2Rhlgm9wp/8bPzPlPuMI034MPcoVhbCvdgQbAqUqroKY6bAjJyM3J5t54wM71F5ESa6
odv83k0WwhsjxvNQQfkuM4rLViNdI26QIiXLIw4T0/EBgx3yRG68Oo39+TEcfnQWXjzLTEmQf5t1
VZnbzV/PWEHly/o5YGrdv069gf9BJy/vhF0ppnp69zfCoQvIc2S6Lr360UjxpY28+ijLNgN+YKma
eZVHLlBkxjwx0GXZzbtkXOpQ/BSb3KNxYxVqYWj2qz2qRd3yUuA21MLbOTZjvTKWGRDUd/0qqTts
6R8xYlzFSX2UVzTlv9mL25UXYkg9bzHoTcCrYf3ejSrdo4CLD+7hTMHS4hWdx+KIIIHX0eJNkLuT
/UzVVILZ7BiwSD6Q6rHG5itJnfIQ4mRh1UKOgn0leYi7seq7hw81tXdABfGlce8c3eBLj8nmGdo+
tKd3I/K1rXmHWDvzn/IuVcDQGkaCym01KNjH0/QLg+j3X9Q17KPwja08O8OcpZVRTk2mIyEFVmJM
DJDtyUyLZfcW8dW70lIQRNR5m3VrKIqdPR/tUwxVdUYGJ0UpCAQxoXiAU2YKjs/ISqXVl4AWmwcf
pvNozZxlvFONuXhDz5hY/ZBIw+r5waFPTU2XG4PiW8upiP2qDCXiRGYH+7Yt75i233xPHpkPKx4L
SRw1hCoCJRRQe6UfZtKCwAbqc205Gf3pVFF7IT0GDFOUpkXCMhbipZoNm2/7oh3ymkreE8YbMKBq
2ILSnw/ILWOHBdNZuHub4gAK1Nh/rRV5WwNNAzE53/BMFHz9NL11MM4UudCfKfBJqNEZNO/LTwTo
+TEqSWapsZod4CMFZJbRBw+PJWjxQzntZyOFvlCCNubF7yGjtn5ymD9hCQnenZKmBoEDf8WhpQJ4
3GolV/IYlUQZJ6H7tevr7cIitFHKgC/xMUzmXdNXK0B/kPexjKzErixJZ84c7wD4zKiWnTUzaf28
x0nBs0cgAoNd6dWlrVLnTRsxKV216Zw2suiyzokfzn3S+MEk5dplusLewJTJ1tkVcdbsy9dJyRWD
B1Ne/FtkoE2USuiV4ErMGoo/drTD+yOwSePDeXFfuA7buB6/JgCqdbg6dJFgMb3NYr8CrBVBmE/v
Ik/BEoEfXw1t1OFdzfnscrjJnPb9VBVFk/nEb6hsuKFqqX9dDH0VKQDzPIO3gdK4HaKHEhCwAx94
7+A3qYfRgo+8yAL4YUUfYB1EeLMBefPae1+DL93+kml+EF+Ea1CC8RrJcuLqcpCepY4wFHpxg4xh
2Ni0dU9Vj3+th6w9f14JDa56Pdze2LzkavbeZuadgyiptL90rO71efFcJH5wovox3UcVVniuvqaJ
BaD5l1T2NN5nqlllxs41jpt1dBAZrTmWjqbzx8TmgtB3n8l9pCZg/yA170ejldFvfv79LjJBt95K
7ZkYkAhEfMHM5XBnETBuTAs9HsnYSJhXouhqI0XlyHY3alcHZOJkbT9H9T8o4hUj4+0zD1NKyuJC
eogI2OqKnvTT7zS/6ruBXgGG2VQIdylTsQtJhJFRgXINCWnF1YxfKxJZgHDHSzDZ6RQOJ53k6XoZ
lhx+SHcb440IKU1j8qTwyZT/8JDY8C4MsnCW00dW3JVQUlyVQxF/oAjQjhPIoHkCpfn6ltanGW1N
BaGyDgOsKVFqRsx383Li6U/qy9XPWEqF18p+eoro5HqbLOg3iEaYD/eqMB4aTgmprBApXpbmZy3M
/Sz3CTbIkyPRp28vC1Qe6YGWzgpICMH/sRzcf5pRIkgzdNPcIUNF4AcbcKwHQALhcQPbnvWZLaKO
NZr9GnZ87H2DQ0Z8moAApqg0nCiUuNhf/riZOUscl5N9+bsBQzoMfYbKgyYitnbFGl4yXbK9HUGt
Y+92IQSeel5VMbtDVV7z//nF9MkaW0dcijnAUna/hAb8FOmI+1ahrfEnEVAQDHtNWt0cZJx2xgUg
zV47HtLT88sbiGJDoVB4Pw1tUD0ArqwEKAmk5dtUrgmubgtQlGuAaCMmnBP5tetBbF2cAa2o949u
4RA7qzutp1WOCtQxzWtCH6eZFEcMf2bb052mSpgtWnT/1B4Fbayt7QZwt9lB6HpDMH84EK7SYpMC
tiJsU2KwT+J5i1rSoZ2NGLNrLknl0w8R7uXUZE9XSd4n6/4YkURlekLtScLezDVqj6BQ+irm9X5Q
NQPRNymEb1J41wbsHC49ok9xGnAoNZIXeqek79MXQ/w2lQVZ6aNgi/qcBxREXXCRuTeRE/xBqrCC
6ru2ylQQfE9QCGAm71eM91UQ0lSX0EcwsSFdqAIYmFyrDboL3aAWJD3w/isEFtOmi/akEhc4YdxA
D2c+0fperBiOt+rM0SZQdGyCCUdzXGuDHPpI5KvA7Sqq8y7a3nY+obQNqu7pgvmQM42+M2PPBebh
zc/2/4QRGmAXarla4xoJjgbSBSywOuT4O3r+reYJUJF7AWwD5xtC3s6prhMIAzAh8ER7mD69Yarm
GXepxaQmVIsRPG8aGA2L6eXNQ8FfDwS6LvLn4gQu0AQSj2rxg5iwfD81x4JgdmvpAbh9Fe+cM195
AS1uBP7T5RznJ4Zd0UTYVQCRat9H6zp8dMhDwOLS54wnmFQ0AeSGteBVI4MS4ewkkE+66uXDyEWN
owl2hs/b9GsyZJzraLJiFnlYTTb0/RO2JhlJEjPBoezb7+6O1UiLzmgHmUA75wzTePjbrrrcfAw/
iCkTzVpQW1C4WDaWMXPqkxIjf8nJfTM0O8Dq+6JnoPLeffr5OXJx423jUHfAhDD26tVm1KwQmb3V
oq/1rs7M/8TA0Y4aU7DWwfRBqwtsNHe6GWooMKoxCRthmHVNI9+flI+33Pjfuqu9V70l46qK2P9P
3g1GpWgIB8p9xliyS0k2092HZbUWQeJMvyZXoHuJrEEIIpSUy5NNx5wAGIqqUolR6moNDh45gbEO
kGlIaUwLq7/wpDLpsjKhE5n+9SkSi5PazeioJ5/hMNje0BKXf6gat+gx+jXKqcxTLPZJ6XF71yti
kS06qD8K4aQruJKOM5VWyu8wvLlTf0sAvNj6zn/xoo7I027DGLb1ReEMa65XZnRTLMHLvRmQ3yV+
qFh0e1tzkK5QM63JIZoA12x7MQbCYgXEsuhMdgb8u/5AX6AOFPHDG+a2Uv+3UouvLz17uOuMGxoE
GZ2vQ9s9XA+K4eMG2hrG7GmGUQXB34pCEzNnL/ZEGtnwfh6vd3SyK1BodSnfTisSM4x6ZZHx46Hu
ZAdwsBiVgEEWtE5uJHM1ZhbShZI9Rg3X+FmazExYqyMvucmuGIiIMNf37JOe0JLSwFWteCzAUETH
Df78ECOJsXDgune6NJSj56TxZG/c2tB7Q9VJCSKYJ4p28FU+U0fH6G0rNO5IKLHaKOvAdTv9fNAj
HvW423T6J+VnQUC21cOF246kUfRAK/ziLyL4Ub+25qhPo1HozVFc4YnbLUwMTewi1vJP6oSmMCbx
Jk297oZS2AnH8/mMeZbGEsE0YaL2F0jgqzP5alhfiVsDRbc2EngHuJ4OdSwkRAqBn2pSAWJRE8W6
TeUrZFAWE8/by3z34HN3mfR24DZx6DGDm0vHAOPtzh0IbmAs/zt3AdkJ3fEcRVE39u/7vfnaM1FZ
Yo+i2eEoa6NKG3HUy1HtniOdDeL1m/AKKKS8B1pZXKdYxPMaM3YWECd0BfUJRJTUf6gKxAwLHc7A
2t9FSRyFDsKXYOXK6GI7sTxup/7rBYh7VSj1DYvs31TDChBK7Eft8lyQE96JnRLK2zJII56OrHba
gvtkvirOii0fZ+Nai0pLZIqnsvy/vxEV1rKTQu3JcRtbBeb3ZuswnpKR+pJKItjrq287X26aZ/gu
IOXADjcvSgolggWc5AdQ8iqxEX8ZGGKpibZLWr2g3EMZBQXp5tebK1VjAW98ysp+BZQZ9eZ0JjeX
N3y5u76EEnjRp1utCAI5T9QqF2c6hgcZnUEmOTFCxZfBiXWvUQfCumEmLLBit9A+Oy191es4mXAw
6zjuQLr3erQMffpPSLcRc8VY1Q0croZqlW0TA2hkwzsHCiFqFhP8S099VPrCyW3RimpGMJJjyod5
JeskkZ7Oqguf9H3q5EOYMEHR4fO/GYUvvCX1uNMgQvHAVWHsRhSALq5+1h8XwvUfSUZKUarlzSnf
JLGi3+ewhQ2hwQlKB9IPgZpSeiba7Z/j4iIrwnnw6xGtx6l6AMi0WnFBQXisu3Wx2ArDsFXBFKkz
tkUK4alo5VDZ5mkasNODv3HQS5HiOhFxe7O+FL8BBzNgOP0mxDuM+pBBGp15nH1tx5uNrwV2zRT5
oyV/GUjBXd1XnpJSs2berJQJf0hcBjJ4B5oU0HN/mpI+ZQsZosYiH52ru2/FCnKLxfBpHKtoNAHI
Rh9942Gs/KYd0q4FH2HQR5lTwKBtuCgXhbO/sEzsDHL1BTWBzULzGQL/p3Iatbg1RnAbcnJqdYpl
Q8HGhNHrVwAKr1NFEyk8nml+vkbGHHkpi4+KuTu96HX7M9zGKfBzUwh6evjSw/ivM71u6G2M6OIm
gMAEZp2gEySOgj+J3cBe//cXJvHa20QK8Bv0uR0i1uvHOfvdTx9kdWxJyl4lET/LmXGGdhv3xXy0
/5XYnGiCo9gXng9JtgRFiwpwrxFUJvRbG6ymabYWqMLHS9bM3jPCJHIEpm/L2bYrPAmv18C5ntiI
sJqMWPCRnUZxnd6AJtU6y1lQeJBexGHNwilO7RlkRdwuS1QeExZb+61w3e3Iq5quLPfNrvnuJ0s1
Stm3dbpLthFLle2rLNrTjGc6/RQJBfjdP5kd1IKCqx0Hg2+uOstc6+y+Tcd1d/bCKTwAbPD2goao
yU+k2kCR4f/trKYhiCTHmNzKvGgKGoQmIvcLpF+U24smOsABD02cwdJiDART8HCohr0Cs+XtnzUd
SFe5BQLbrEQ8gjTsjKp4nkEVA5ScSc5N/I7qjOIR6PUOSgRVfREA9HYIlZJrUKZysT4+uVPvdmwJ
n3xUtqzr6uPSSDR1uSFnmhJSR1nfUmiMxLpi4d9UlgMWH0OzbN8xJ888nzoGQau70rB8I4VcbLUF
ikku7KE2ATPR5UNFegoXWxqCxnag5as281IH6c6o1L3hOs2GPI8dj0KFxiUU4Kvuog/MUNcA42hO
+CLadKtxWR+cdNIsD/UtPT39wcsR9BQxXgTezTSSwYmp6O7rzXH1ykCbGC+umtrgbFDcfiNIretf
ouiKMa9waEH51T8saD0NM9OjzELYy61koInQM3ENmdeSPqLQI0gve4rYoG2+5rXEpk68gAPkYJ8G
nGb88RjN5jmDjTvm3p91Hx+iBiBzEhm7Fc1JSeB50hOus9qEL//wFEo2v5HCKdns35hEujJPqFGK
QGQc5MdVN0AS6P4V+a/dR+zqKEcr0k7dsF5YMIofGvf+z+QM9+vqvCLVz+DXSBwN2VOMc7jZcf/u
OaJBJeHnpY4DKC6e2F8ihk+OLmzBT5OVKC3RQxQoBiH70m83wgYDypScdDNpRZgnWXsKnwOr9OK+
lezYZvUXG+rHeKxXbXz5OnMYBYz4Rm58UHJwQNicw5d3cJD4JBJGQEnBogesAJ3GhBoUiWTfOdmJ
CKn69gRhow4R7oxbIe4FDrJyV/OvuEXnbEW4o+Pw2B1NkylUlMBi2lihBzdY8RIm8wEUIS8M/Uqr
nFyhFWwEJu83lxG5ourswxF+k1TJAvNigBeZLDGfLISG3WMXcljE4jXvhaL6MDu3blQGb5GDUhpQ
cx+8qxUmdNEf6HOwh8A5tV/47xTyXAPb3LF+KnymwuvD8/IVCW8NC1W+Kv02pePe8Gag5Jv4q1Gj
rOEH8WpgOGz9NqynyoiuF5xObrYwBUKAiaI4kSwSOgmUSy0R69UUK9tUtdG6J9/8gSCr9uj1hKJR
ZIh+InGpF2AC+Usi7CZeg6fpM2X9PwCn0Y/gW2MV0lc69Mcyqxu3tppYPqXfm/+VF5FWs2noZe2l
6AYFhTf2vgGiPKUDGe02j6u+QLSz2yCwsbfOjktYcF3Ie660576jGTfzw/d78HUmy44b81wehUX/
2p1N2kMoTYpmzZbWTavYtS1iqrbxqwGGGQBmK8+tvhb6QQR4Hhvk9FokxQRuU4owlxdi6YkYVEi6
//iRNLTcszxLo25lkmUXM1iLAqx9bh/nCgJhrUR3ZAeWITo+AmsX6lJrmImrn8wyKvNX1qpe4UyT
kZksGVSI/5vJkiFsbSMxrz3pBh6bn/sbFe4LjF0yYRQv4N+odqwI9Kx5hYdWSfyShRM7WaJMtszH
jFpsdUTdFrXBlO1oSN5phUXs+6ShsNsX9kZFUhMBTjAMJTZUdrFtnJJFiA2bHeJJMyiozcWNonfL
+1sjx4pELBclXspgTm1YPXlTM0laDp2obPAWXOAPGVndr0TFlVzn8QB/oWQKO6NijVMQsoYix7ST
1fmUf75G00/f8dyIj8RFTNlvG0/meXrmCl7b9QaNBIaBS6t7eS3bwNCTfkT3ICFWeX59FFnqPh9D
3LvF6QJWjvYnIYr0/ju9c4llFBqiJ383ok9Ay6YwQfjMHnxqSVREhyge70pZ7rjMB+mXGffAUc1R
pPYdu6MGTt18gYCHKYGBzM5OXs1Nw/GkC/24sNeVmwnpXkpF/DIbj3Cc3SMdTE1FMTSKFKFrv7Ni
0KTbvZF/QGPE5IlN4V/UdSQORKdsdafPXVtz4aNxpQZ3qQUMqWhX/1/Cr/I7VexVBwwmHvr8kAwc
mtgnEPROoDkkq2QkqoxUA67TrF9R92rfiSDMI1rkOcAra9/wcBHJI3lPx2EwJDB63z+6+nTgyxgz
M0I5tGBp6uj/3ujzT/4DRd9qs/3sOkCIqwXT7+zYXf/Aj6C2kvsmxD13yedQSDKnPAbTCmnWQN0N
Q2ffgV48XToBW1XIgvviC01HWhdSprkrVnxLFN3h0wnjnDc09Vyk4DsaJiYqFs1eRU2ngMSY2DSE
qQYopK/z0PaH8EVCt1T/WV9QRC7tKISxiDNw6ko2R2uDJJGEg9XDpsbj6rVdAd4RmgtitunAvTR5
OqOQrifWm+U9IEJ4pHi7QggzOzrR73qs/+/TL8FXhkny6kknpTArpj4pGoCGn6I/jIFiVY0VhdZa
Lfw2IZUyHvx2URvzLgbBV9X+wgW0F4/kgT48SdyN25hSbfv04xrBayO8y355STI5qlaSPeYEP6fH
iK/FaAarXHJywsg/jCsvM5WcUTjWW1lczjt5yxYjGgM6rfYU5LHej+97w+2O2rJ/cuG+ibrU9fTo
Re/WRVr4ilm0pbP9npLZYJ9BV69XkQv/y/BC8LHf1NzOqohFIHGnjspIXkny1oys06U83OIT754k
dy6RihssIVb+XAiCNRXJW53yFLe4Fj4gNhcmB0a1apJlosP3HtK/Xk1yb6cUjXJwyQ9uUn+4aw+r
hFeBzTAD8W7+ijXImCiqStCo/1HRR14o1J1w/qyQjHsGioiGqkm6zyGd+xMt7+utlJ9WdMrmSK/n
TXn6sCRdVTibFiczu2JdP3gelQ+oj92qN5rVub7wtm/lae4CWDFr0Ea59fpJs2t0jAmXnU6uqdTb
E5iFAg7ahLslWrrq7JOI9LRbZRxDCHegzs+AYrch0GrWBIh7pubjkQ7ADumJasYfvGceFoC+bTGd
3HWpzJasGcUWiUx32BjUiDxmu2m1CDHlIqgrt7DZI7LqBzTclRViElxGFxrF/ol/ZX+3zeaQAqPM
S1Uz8VjFqE2of6oD3/1tjE+k7D3SsSQPTmFwAhc0BowtjFOld9xbfyZ9gmZLZtsxTlsFqnpNWe8K
6TwCQd4iscXMxNj8UorSyqkzsfJ/8FMqqjj2THW/WBjib48RWXQKTAoNo+zxS5wMgv9zeGy2Nz6q
ZknjtPOAYLNdXXxxB5QUYte2trbsQYanClxjSb9NHSTMbc/VWPr3FxCMofsy/egLRx3bZn3gh90W
VXH8GUwoWym+8fGEN4inwRXImrLaZIRwSpgUm3YERQ6BHA7cuPJW6bxMvitHLcD7VasE7GvrPYa0
faeAix4QfWgka7Zac6PqvYS8OQQVLnux65pDcG+cxRAvrC/F6bQMoHt32KlclKU1aQBJ5krh6szy
tiszOtSSc2yCrBZmgsRHhUbGXJ3JPstopcPELfIHbmnXNoHSXIOQ7KPEFqVh8DpWb9xHeDBFst/G
9O+n2wsoNemVHIo82G4AbCsqcdm7xzLMpnfETKlscxB6FEgrWTR+2HMOFgb1N3As9Hlpnzp9Xtyj
dEVOOU4GMuLYPOtc0SYvXbNCxMQQ/qxrUjDq7dA/fjrRjPpl5BsBWakJX2eYH9FkcdBxFRStcU00
DXHeLsXQ/8DLXEvHSRUBSF7xBpNUQeqE8w+Btw6p3+JuPDcQjGIHLUzveIRJh84h9XfKn44YvJcU
lI5hn3zl8xQSmBJFSHoG4dMBXD/2mAQuzBAjS+cZyj3GBqhv30d6Ym9OHJwdTQFiJWs7mUzmow9K
1OPOshgWQs7ITkmF6c98aOEJcaMX19wXPlhocQsSJIUDtwiFNZCOltgMCP5QrYLcQy6+cFgd1Kif
fwfrV2MN/oQbxkggt7m1RRQYsOi2SJNah6YndWQ0XVSw7o31RGOVtke27NvttF2Fd5E3/xzLrOxp
g+WWH6c1CwTQIWeB+IbqHXUNMQvba+3GFkJKOfMQ0MJ56MbI39foq/14mFeX+DCe/U7kgKA7+vsj
x03/894iOA9D6g8lGnIPE8k/2Jo1QIvUBf2j9ZWAANRD0mBekJOcNN6Z+B2M+4gsr8t08xVSIzEj
mPfCeX2H0Q2Apu/nHM5lYJ6wBy4BtMbc5yy+ZLHvTFkTiQRoToa6K/rJbwCA2NZr4m4BwqF8kUWl
x6wREUJwfX++dRR7yAdRAdDsCUDMGO3mMCj/VikJ2He1Jb6zV28jcDMNJbI+zMmcVhkfKxcWIq0t
l2abs8vDH+Cd168xAJRbhsRWYY85woD75b1ITNQRdYGMl7iS+K13iGHRW4L8+AVDAkWERtjRWAAO
Jn/KGNs0+AUXVourwGFX9yH10Zxy6vXRK8vKo9+4kc2GhS/WJUc17NaM8qq0+7G7AkJR8qq++L4g
7g9y5XLS5P5ldlL7jktZfmAy+0PxJL3p+QOeikBWrpcVqkAavtKRs+RD9+/M5qc+X+VKDVJa2Epi
Wwr6HhFDhzCCE2D6Tdt3MSmwo7oklyUc1JEu/lChonS+j3Ae9FaJJEdc4Gg8LN8x+4fyJgQg2gvR
JpRUw1jvmVXt22fyxywgyUihbv9V1WBB4K57bEa1GYknte/RKMK/C1p1iMhyQgTyXyq1Bf3Aj7+I
7BS/vFPHF+psWXDUG90BYGhcdhx8FRCNNOO+34zXQgVYOly9FlvzBpnsX0bTk6vZrGpk51RWDQQN
2c8DSy+44el2v3B/oPUfPiZFT5lFN+OrzBZo+vgc/ba9Z/ONkclHMCbeFiDu76Y/VvqpHgCba/MY
c6THoctxUDZGTtnvzA/Bynj53rpXZ71IeqF0TsVVSQrL0dvw2Vxjt3HXsKYAq/gDZdjYvpXeb50V
YBMJ1+76OOQhW1IYqxyiXV4nmgIQHBhUcc+MRrcIv+p7CrunpWfoaQrDJhPILTkw9zvu+WSafh9Z
KWBRKamcZFWgKc/L34mqg1KVJ3Ey/+rEBXncVvD3fIk7aqZ+4q4m/hgae8stgXkY/+mzlc6aBLyG
Cm2NUnMZqMfpapF969BoMObO0W4r0a/gMGNnw+7o7IzG8UTblT7S7ecYSdd6gGr3aGSmRa9X0MuH
WCupPT9oG/vVlLo5WD/qQ4SEHQctL4z56O726zdDNNhY8WLl64Mc+MJw/U3B4SZdN7LiiUGKd56A
73kpEut/7g4x39U2m4vh8+aVN4cj/npq80tCtsWqVymVcoohjoEhKDNNt0U+VpVOZ9GOflbLAbxE
sQlOTfdp72kflEnGTBh34atTV0VI2K01y5rH/ONKasby8e7OsQ03YuGBnNRnTS16w96C8bkEfqTS
9ELdMQjJV3qjGURQZV1oU+lRyudc2vQ/Zkv8stpI78twyKWXmErH6TOV865B2Z6VauxUcwsiQOe+
ViSpE3yajOmhE5wT1s/veq0oTXI3FzB78KQxc10VFKZeSlMdU/kVKkhwRfUWREPe0OqYhJZN3iu5
xZc7NnPAkVk0CrHh5ENQbpcC4b2edlqU9pxIWTZfYkHxn8+LFYOcDNkPkaMdm18p6SGkTnoC8ojC
pdhZEdh+M++zkWyV0VTN+NACtI26xbL4ciIDdl4D4yhiKUbn2hLWfziQsWrQ/j3z+hxaaJEazc9B
wClhERWFK5t6EeGLSoxI5s6D1jQBbg0UXznmHqi60o9L0w/60NMlkGw0e2ZXb94Z8Byu5Zy0/mRn
kshdaN69NOCHPXMeN/EmTrhp9lcW+2bL9Ym6NhPNNXu0UmsqClLwDAaDQSjye9kD5ZnDEMGqz9Oo
gcMRbgu0BH2vs3aagXF9vCuak9qB/Koe3FhrgnubXChwlN8Wz650LrHCUcU9wo/goltYe9wR9iT3
NKT0dH29nEBdgqMu0jO8DcIO4X1BxfVri4JziNuWJbDt+NxAHzf41H68jbMcc+uh2vFtEdvKokEv
u7+Qw2QvFJhvwieEnVsxh6ZSrzvdrbU2m7658LqzwavhmBPHaV/spSo4do+4uW3BXy6yH4d6lgF4
XLLxIRuCqqpo59NbEZ/b+Xq7f6dU6oz3vEnB3wI96P3VP/Z2QIdpXabO4+SGaDqXubBJkX8gg+zu
NgkK63DVWq9yw7xWwbQ9hXybgJkzfn+P2SBfJLkqpDhzzwgJnCj8RoiZdaX4UTTBFzmBsffKbCr0
RZeRrsvAeg31B3cC75HBDL730WKjNoTSLxs0cIrmK6zTkP2fejnT5KsehCg3nYGGHGrhhZRHgjSM
ssskTDg/rcRHmaYI49z1ZHw/r5xqOfVCjefgVKB5ZId5k1vtg3UHWzk5zfL4ZpTi26FSC9a941Jr
F8mSAHrRdIp4t1fzLT4M0VA0w849lAku0woI1tY4lpVmnVN/SouC5uAyuvbtaMO6vGT85qQtP1Qa
zicG1Q62zUTjXzsV2fQz1elmuMlxAAf4d36oeOZ+9USRG6TsG0iJzRyCvH9HA6wbfc153ySNG3zi
vaboLLpV5SYEWaUsi7sPqh/Zwn5Qh0ik3g9k0nhxoD4SU5Lb5rVi/u+eYkfj3Q5DRvJViFGJfeuz
EwFqcE9wc2v6e6qEBhQ9KQ3RkQMXZaKjyNAQcvpegULVmdQHSNuMouOaaRY95lxH0r7D2NLt7F61
AYMRomV+OI1XQ9LhjsdAMg687FOP8OGPo7wx8oppEXZ8Qrd/f7wCHMYPnhwgEkEV5W+1VzxxkC0q
Uj+resLS5YJvjj4kbmfEH9GVPilvU2nBZkTtayu1eKSYWWW+hhOlK8AE515pB0Hd+vgqHZ51Mz9g
N1djC2p0S1ewJRsEBcarCpSpJHd2U/lmaD4sLrOCau3DIR7l42CT83CJUkaXW5w313Q2qtkwrIY0
b5aZkQfTm8JF+5PDB1NDjwNbbcapMXWz5Rz5OxGcbr3Rwo2nPmTLFxqW4Ft/1gi4dLHWa7UnCVe5
dBdDxN/pL7Vj+inYa9mGhJmxtCrUWh8jVxDErFHDqt9nPy1Uic/i08tw96TotxrCxaOnJizjd7Ir
2gf7J5GWo4xds9Vjkm58RvstFUx+Pld1Rp0CDZfWB9prhfzuXvUl/itxxYNbI1GjI9c4ho4x8uF+
T7BGcTZklR3GzUbhzPHghIP0GyUoPg4r6xPOoJ5Xjd6/XnEaoP8tpq7piEVvuN7BDW4Y+QCwhDue
TrGgEf1+UEbHDPgGxfd2Jj7mEHVsX/tpCIuJTxVVz6ypJVr2LZmYSutmfxgHmhXL4iYgmiMSCNug
IU8HE3ebKlcAd14fR/R116rIrYJvkpEfhK8Nl4f+i3/s7rXC6bh9GbSdwVRN53e/vlUKEzW2GR31
xgWHhmcKh795GFgCIl8b+vB9XU2V8VA5UImAKcrQVq7Uufh9962iEq8RdWVndeTiFNhdZR/rhAW4
pIhYR4KgZZzWWmuuBDTwTOcD18Pyj9JRFA/FwVNH7tCbHbG6wYp0a0uEiJb1fYBdrC0ymmYphBqM
VkWbFGH5rkfByFQVHnC/NRJbTw9nRtbTB9TLXVBaCcq/edHtXi5CZNDR8qdmLvANWNZB3Yke9uDj
nftkETWnLfZ9/TWz8Je1+p9KIFgk9LLAJ4BrldxrdgDnHPq+fKxj6TA1h9PRQxpvpNqX86T2Bqxj
/gqtLqA1MkS00DKG6ezX21FFxLMNpl3CGd4QGs4rGuKItlOw1KKrXsTzcG2Lecaa9xxpiWWZ5FFq
qdXz18GBmUXr4l98eeASS6lpK9qytQIGfp8aQW++XyY/KNcwTsx60yw9meIFuASI9dUXtOcgRlQR
oj89DyE16iScJjuFdk82tUYkuRBWkj3e+9Vp+saMsxS2b9IQ/0fRqNnrCUaOmWw93HQYZXgLKFFB
r9B0VcVOn+qw+VM1dUSnoqrPYCakDq4CUatayWNLaLT4RlffDjer1e0FWThE7FS3rIOOu3qiFg6f
LjJs1b31lR++TyiH33UMdRO13qXLbafvbH5oyi2hur3lnb0Ink+WPdlezYDh/FVzsu9uvh5vT/kf
NQQr9nVD8jWZYD+Kf7MiFFHp3D7zC3jU8lB+4lDM6ofyNhLzTTCe2XXcmf0rjeYFV8z1uj4wUlUJ
YqD0ZXkyERFWtb1BFMLIclR7W8gU9//bsZCgCGOEhlA4JmHGjg9uzcDYFFSaEziFo5SzfJffTbLY
B9F4mEJrkfAKZAiIRbf0FnTFuC2SgT3LCe8ZUdGEuopw1DAkCW8+EnTbrNtyaXA/7nxyHv5rP3Ja
1RxhaqtlvcxgAhgRQ+ar/ThdFivyuex71nhglSyj3BcgBOj5mzGoCUJPGem0BD91qImCUDEnp+w7
yiuBRnZ+w3N14WTD3G1PFzxLMZYm2R8QiDyq3jXQvp3Q1U9ExTogBPiabZSSjbljBke88zOqx66J
eZm/qJ9CfAAcsi4iFNED30Lp2X5j2pvKAlFNLgCCvsh/oo1rW2QlU9AUIsxfjCx2ZE/HhdxfUYjb
TxaNVPqFtk+nLZNfWiCSC5mH7ozZsnX92TgRZZc8Olz6ML4mZYC3pjg9BJCTRJNwHye1b9VH/vfl
0bzXVQ2T3J4iQm1k3SzfUVTz/QrZPXQ+zR37GyUGGARvdZnB1xTVGe0ph0wttG4hLmcFbq6/urTf
K8E7cgWIrQgtU5r/7XPxf/fw5Hb+b0ghVtX0Alr8xmZlWYllhIaJMoO0wKqO0SgVpaTlzThXKMvh
MzCgMKYpGZ4mRNXbhuSLZmm6IFkTeNFkxiP1ne/HRiHhlvnQaRQ5t+NVhGgXF7M4qakAuY+oN225
Wb+NVwOezul6pfb6SzOTTJ/GFdgUmWOjopnUu5TrvqHMVO94exPRNftur1IdMJvEKYFHajqZ7B0P
zmfC7i+fUWN6aWIFpOnqM/JYVLVkdXsBBi8J1XIZGTLzcoloKnMjIIuqu+yQZYmMvzsVtZXZGFwh
O7iAsrWq78Cqel6qC9l3ALIgytVvvc8ylr+Y5BoAZW9L72c3iMJP7o2Ejr7mR9UX0mpqhxzqbtYV
9Z7zK8k6CULdDLpJJfjqX0e0UaCHMjr/UnEFf6pbgF9qIea7pF9h4pe8ztDt5QD5/ItO+nUN0y1e
3GqUm27/GCACW7jK7XwZN4ojSetSMs3feVGLBal972zJCJxZrug02YZiiwQlahZzjyTAppoCpR83
hKA5DkTXS7x8Q/sZkGu/oLtB6kZySf42geXE+USoTaD/M7Y1bOBwjEkjOWq6lMOBdzkqfWNp6nJA
Ahm38j0L/5gqbYNETTqWKWNiovUNiM8mNbh7HkkUiY34Y1WhvOJBfNEfG4z1ILKASF8z2iXrJIim
jRTAJjm3wYFU+ZPm58SvIVcEWBnjUEuTzHcinNuGA9ib7CAYkg9VHUyMg+ZDzu1b8mqtTc80MN+C
0muldOK5irlGkqTSOrfeQfVVVObHpUx2MxnmNDtHx2+xBCYlcuhNNFCWaHpe5sW/vrnM3NVd+HQf
R2thyg+706VRkjRdMMnJhspPytJk4TFp5Tl50WM5bcvvDzoN1Olvr7DVSiuisNTCPxQWM/QuGEx/
ZNwvnSuB/IsnDaBuc5FvyLdwrZujKV9YXUj+xYGLbGAFKqO5w75ukmW/ce0paIJD4PC+LXhjAfRv
dpVCvuzQLZvXTu0bxcvdKqF9C6lHhP+utEMa949+3HaxIaUtyyx8WTP89N0GxDekQwNGR4ezsHxH
Mb2GN5ebljaT08yhx2RjSKfbyENrWe+LyaR7UB2Z12kvQoLpL9JlU72lvWju9kybmzfSEVC6F9KN
PdFpW4N+qCy6kmypc5/GR+3mWJCjDlkzehoWahn2hZ1+iaA8PsZCNkeWZYUAZktSbZQMLNEfhmij
FLIDj8+lWOXQrGA7svfkuS+ercO2Ji4uhgi1+T0abPvwCG9Ev6oCZtqGlr2seD9SGxXXHju4OimL
nFuMR1fD/9wujDCjUYTRYhOck0EX26qfPPi6j1ktqUXYyiYfHr7ZJJYfRUBPfqOiyhubs0pwkBrM
pMp/YMBhYSq1iQ1f0aKC+Z/CrOvIhK48W0OlyQif3VOBh2m5tW64bNF+bV3mEFEpb/3oWO4qt51O
ClTNKsQvzRoui52BDnx4KCBCiSFuoH00t16wWKoraShk2iMd070k6aMZmgapyeiVmMJhfICfck/7
d9pLGqZiPe/tu6t/u62/uqjrIsFQWWwc93mK51/rBHbhfTKiWCcMbzhMC6o20n07f0+wlwN70RCD
uFAGIv8D/CtqDmd0n6arpl9CZ67Go6dhVO3wy1igDRfR22oHONz+8mlIeu8oFKkAg4R2NBz7qV5z
6G7K5M4ZKMEOkBxY7TjE7lrgh8KkM5KEV08Mfxm+mYvHs+vzrW36nDckQOmLMRVFRI7mxSPnTj7s
1kdEIQGkmHRr0BNzTcOwXi9cmDdlHNtc40bwm7PdSf8uX2OJm6YVqNpr5qk0q1thwzL858u57xoX
hP6iqtgpc+nT5ANT7VArcUvhxYAmKLp+zeXKMNHQAng2UMiyqBB8l3gps8cTpxmrajj9rhjQxmOo
xbgZw3T0Me/47Ho/FphfgVpInNHBad3d+K/nEhhkI9ThGewUI90kgPdtegAAL8PqxO29IDVWKD1C
wGTpLHI9CcowBWs997oP2rKSyvxOCGBHW5qcgiOxRAId8Ik60CBNmvNW41GIIOuuHZ0xXsZHfqUj
Pmj2b5Ft8bTY0XnmBlibPNGEWYEShb2ZtMo2pJ8Oasht4iPwLzZNDli/Ev0PHTHGob7FlcSvEDbG
cZNRwLbx4Qy6+v2tH4GCKrfaMRcu37OG8nI/6Fayoc4ie9SCNIwDFQKyvma3La9E2RF4JDCa6/Xt
TSTnAmZaHBw2bf0NPinmHPX1FD6GSWQJ3G/sjxwOKwV7yFlVeLnkto8uVCNiUKCulOfnB2y02WkN
ZiHw2Zga9PHvy838s5QUJE2Iyjjcuz748py9Lla4nsuL2ajHwP1vA94jYxgaQX+jRsSejJRfLZLY
Plk1BPy7UdTaifXb/rnENn7rkLvVBXTn1PCp0EAMimc8tkemApcRh78AmHw+MhynAwlreeuVEvXX
QBq0LWB17gPPe5mgZgTQ1Jn0psiLTA476M/BI0ewdmxZOJr8YhscbrhJydEtrA07aeZns3RVhWnU
i0YVozbRBQgaP6ctObPIGxNyQ10nurxLR+jIDGdernNy6uFoaoYM/Y3fJaHQKmv/CZlRokXoFiVT
t3zJuR/BXKAHvL/4/+Osqjj/8TrU+d6xvX/mQTCwq7R81Sd9+cRrD90gGa4ANjDrHjsfdEgPbpq7
8Q2sDe1P6SfGXwzJcqPg+kPAxe1zdIfU2/vHDNI4Dd/t7xShFPjcXkQLXuMjCclvVtFMoxAeJhZP
RhvFisVdv2s5G4uh7nfbUDKK0A6uzo54/NmQTnJAHW8k5aIl9znYTrSXFEv8XEw0/HQDAO+Y5WLw
1EK2C1DET8IV1NwfGg9N+tezwPP59cmHCXRsrkJbso60es3v5/sU8Wp1fd/O6FC7i3uDEyV1+tfm
UM1OfdjTiY+ce+imn6JIbO5mw73m77DA/JcySdsxEt0Uw0NR5hptaclJSp3FuW7xv7ksHuLg6tn5
tbeV03x2elz3r6ZPYTFzMkySFpkwcVHx2pYI2izQb0qi+ERKggUcI9E3J2Q/iPlZlWcJAVeGkuzL
9BGChLn00z1QhSxEmj48K+miWmQxJJNtNga3rT5gyyAgJkobNYmJUGcztsUYQGTqCfwPeB3mw/Pc
YKInziQ31zd6yfhTa2UQGjdlNq+oWWCLShSd9skxxRgMCCm1aLDv/Fplv2S0mWKysdO+XQkjgZBC
gKSvQQmlDz546A+R97Y2b8HSUMIABsxWlXTdAXLCGXV7VwsMPDTbw+crOSx01Pypv8vQ+pWIlDPq
hhwn9YcLj1r6MVIxztEhIJXJYawjV8S0/rXdxFABj0dg9TFanapbgCtSmAknbxrX6Wd2bnDxM5m+
StGVvb0O/wYZDzPonwAa+q1SpvVhkguuqNPV8C7iAFbo9od4TcQ4QFI4j1845CZRDCBLZJHcPMpA
QTVu1cCrsnnBH/IMWO1lht5O50FAIoxP/q0jjKCl95IjzDNy4FvZCpgs0yknStO47k1TzB6LZMFg
DE6PUDRU8fetZcINVvXxNLb5TiRn4u1sHTlR5QVIdlZDm/AivZQHifQi5b533NiQpRV+nc9St/aW
slIyQ3p702Kd45GpfKc5EeYqNfPXl5XhQDeOX759agOCtwTosx/avI8RqqyDs09jAcDrAAD01PvY
pwVrF8b6HXQk8NXWGdwwhVFj1c56h50liIthog39JKBcnNcnKYW7v2avGkW4aS04RUCPPGzIZxgD
6bV0lYQ5jnAU8kOxEUcU5aWkVLnS5B1QgO1mgsI2vfKSPsCW6mgggf3IHl2lkWZhaEpxapSZnmBz
UOAyzWrKDZl0eJvoScg7uevE8JIlN89wRvmbGAshVQql2p7xrfnkSYqHnUUDD+kByV5iKEVVk1Qq
LIdrpabwbtp2ZLvk7hYPOxtqK65A2miymQp/hOwBHKPW3sGTvTbXBuTryAbLPzz0Je3zHAHUuMo9
atVqJlL8YPwCO+cMx9/K05aTM8IbKpUX3sdEIVzR9Sqbch3OnrcmaLJ6p2GtwVoyGKg58DAcEX1H
Bptg9sOjBBBlUd16FAH2fR72c5l7PNtqAvVC/LNJ8G2Wj0gLKrWusHz90oliZpdbBk02rE2C1afp
2oWB848tUko0EzCqcWqB7mP3xaZMB5Vi/WK8nB3OpuD4MxziB0H94JCV6/bKdwblOcLShpKr2saX
aVH4H0gJxZBg2LFdXWyY+8AJ5PAc328PtqOzvpSACD5oJsL6NtZSVrUfOxd5fn4FAivihXvLqqi6
5DR5Bxvf3o9d4XbGPAZ205qC/W7xSl7M472dQbQdNlOwpPYYd3HXKVIPBwcNgmD37ZgB1H5pvKh5
J6bEWv0D5Jw2TwW2OS9ET17PuMUNjkGEpURtJYW9gxPVoq3qgCosF1g6/XGo+veWAi1A5eT67YJl
4iW4SKEwkHkzqN1Qxes1paRhlZhftrJoTH7v/0EIHfJfVwHxWEuNTWh1ZichoKboWvYYJaIxD4CQ
CpMm7l57ZISt6WOxR1OeYmS4VimuFADPllQg8/fZGgHlO3UIhgq/nc+fHY+b6N9mcLhvig5tlsCl
P7FQ/nDEn354QzCAAEYeR9Le7AP1XwiXVmOEF/4AP1nRfr0VOQS0ocv9UzVWptaiiQQclNSqONeY
HapJsm1pLBQgmxCTzNUESJgjKEGRqiasiWAlzBrdtQPmcXz59wuFNVnvgYKEACaClxCMSDGyipa1
RUjQo+eHyk6cFebaIFv5tMJ193+0Bh5Gv2tSXm3KppDFB/dXnlShlbtTxFYqXPwy/B9Ma/Aay8ZT
lYrVVSadIB6UXowwTi3PR7thVUio78wi7FxOXdQ2i4JqhaAyTYVuLH6KuTo2F7J/ka7wc3E6065/
ccZAscsVfyEnzOGzdLca7t+YM2+wzWhSqTss0Lnv2k3LRo9K/tRZ4vFMTZvJtY9PqR6n6yvl6iqt
c4u4SNIkibmTnjz9XHJVZbnJbAaAm9j4UGlYMBlbDRsLPOv//I7YffoI25WpA6JsKizJgyYMa5Ww
eDuZG/4i2uiHe9Ec6stJxANJIrBIz6odXxbZbDOH+0Y/ne7N5k81MBnTm+30ZwAoWInerKzZV+qT
wWV72fQSwJ99UeXQ97APY6qNhghlIKsU08rdYkBX6cmH3ddSsVLrH6TpU4P35aqIOAhRzPVvWMcK
YB6oK97vgDUxO3mxlGlxFVegqd3dOEXubrBG5WOBBvRPFCe1PPoBm7FCbPD7l6Xxx3xX7mctOmK2
1FO/cQflz3M2LtA758rijFz7YHntfpZHg8in4T1I6zjSKWBuWRkyb4ld0TbvDI3nKZ/x8GrdJB5W
mMVdH+mlefyrYv4cssEcPjFpCazsAX45XY3uQ1/ILteLVrWt4go1z6IqYSb5OgPXtSxMT5eJiUgG
eXON4BYNd9ioSQP5/lTZ4hg6bjJJG0koaAQ2GOUwXilDPLeBfiq6qLiYzKrNtnwQKj29ojicAWVY
4BmyzSShplrTYyantJ3bDmBGeTuTDeX9L6VdAW9UT6FwbtDX/m5S4hzBafngBWct9459kPn4Cb40
9ua33MpnR9mXyYgEJqUUtq1NleG4ndDNoWqj0wKEvhEAyZ8hBFlr4Kc6NN78o/sPHhiBbU6XSnFC
Sdrd73Hpp5uAu8+0j3fZhiDmhL8mXnYQxh8un/f6oAzGOTtlWsLAqZbS9VXGNSMrqKn51TcicbYv
6uPo2QZt+wmHyWf2UlPo3BWa4wl53fQ0sFj0OgV9Z1Ol0sONhTOhPZILf46XbStIXPYP8u8INxXT
LqFniIPD9/UjCfAZoIXPtXIpMaGT4mkqDLcixMvvHkgEb9SiIoJM3uRYkPehH13b4kZofeoymHam
8Y2wNacwOfzI9hs63dy3IJoY0W25BNAAuBjr9Oag6h7JcsIK+0iQXI2CoAUQHTAePVuLg7uMADWl
Yb+65VSQcZ5J+i6UzC+XCiZVOe/V5vA7xMUz8ilzzd0wohMxuyUhU29DDHpBONbf5LpOz9JknKkO
T3r4yiV0jkDefYl2wwkFBLADW6x5DZXLiJWpnXtLwwX6jCmhfEEX/uTYxrRbNitDxIFaIj1hx/Qb
oCGB+dpswdWnQ+T2XdXra8/Dt5w6nfh07mCa9uFe1XaSN4xONATjSNBntXy3PcKdCqjKiRWAMjbN
Q+x9dXawC595lkCFMNovPjtH+e9IwsHsk8uvK6shr7T/umo4tYDnBlNOnaMUbYVZ8PqNZ6gyPjvR
K4X0zuCBIcx/g1FEREZDyNYWIsUvXasQ+KAq89VZAY2o1kCoxaYG51JZhxfiX3kpJB7yYzKXOHPj
zb1/xl/P05kA1e48LaIK1oQCgIe505QVs54tJf0HDNhiP+9si5PYXcvtF6F7zIrr7ijjBkCRBy23
2WnzPHzMFXMEPOAoKIg2O1SueUdT+Em3Qqh8ToOasooUgpuz2nSD9uIesxRqiNljAy6ffHoj9Sbr
Vgq7kl6XcON4Acpm+f1Qv7BECJsIcWe/FSeVuRqSIhcFDA5QSfpzIvKfyzj2XX/i0OHubeYQ/k+C
9vr0vF+AswfTsAKICgbRLZKrfNSAKqW7I+k6Ss0qBgod9boJ+vy293D7PAwV74m3favcPIqKbjR7
8dpBZBBQF6VsoBGxrNkxmZDucLHv2EDnexNdC7H2llbOXsmvkgbt+/Y6j5A5dW5uuRIXNzLa4xaM
T9HQAzmY1CFD5tuYMcEBEFSDFx91l8C5Y0j5mLnEqtX+ne4t51nWAekCSAP4UXpI6bbwWPJeGP5E
MCvQM68IEjQSxr7cncdoS4AKNAHb5+ReMmSJGcRjh9y6N4lysZ1qFmI3YqR/cLsXyL0T1+Flhd/R
7zBToO959RjnhXNRzCWEWSOdOEzpF9pFMWlUKvqo9LS8pjLsdEVl+BVnoFqKdCVHRuDanKh5RF8i
B11xCfrCu2Sg2XVBUFWmbE/KhiiE33FrUn8P/qzb3QTTrswg6Hb+qJnVWi5HZTJXTea23aZqwKVA
qNdpNapHGNtFTVCgvAwDMjgWQkWS/Ifrc/S8U+7U/oiw8S/lPJyYVs/0N3IUj8iDXNkuwv62ilTS
3SdI5Vcm8jiVRq+NbGqHl02DHu1H8g9DrhGRPEBef1TShAQcMYlpjMTVnnI4q/iYSFbcv7edP1UE
MjfhwcbuKoCx15NgWI03S6XYrsUjP4l1yUp16/wvG9sGAbI1Tfab/bCvsw7eZjMucFahGB4g5no8
R+9k3qa9RuPWamBR4CiT32oXJ+Ueu7osur8oEqRagLD1p64UleOy/Vyhk2Eqc/FtJTDMs9M2UyPO
2IO4d6ahUX8UGXr81BnwBedA5LSMk8jRBXe5V1UpOlbuEng0sOKnu9ZVthz3W8PMYyS4ZLC5bxGL
bYcnQqLOEMX2rqhMB247/Sv7iJn4FA38G8KNGwmtrqry7CXYOxop/mKR0BxU1ZIOCSzj1McaNsQW
SAsiv2Q7+IU+hNmoCO767rEM48ENTPEBRp3HBB51NDNYAzPnPrBqal/OCHfba87e7DdOGD1HDoBR
Li/f2LeIOzmQMnI3ZnK8lkXifeRTxjLZRsIVvvS34O5N2I73DAURk5GvQwns8GhITAPbEuHLYTor
bdm5mPDm74OIpit0uNFQzVexLrgebbtBdZFd+o9/By4xcgG4vdLwccWDpkgisHO9EYTHEPDZYdWW
YxCUlEF7bDT+dj+hf7BLqCAFkJIj1TBctN/CrzkHjOkDqPdu0lsl7UXT0c6THDbfP2N52KXMPwJk
AbQl+WGM3AKQa/x+WqtxU/veY1dhnBbUWstGzwx0DwMvWAti3S7WbzWG+/xIAJhxeULWe1X10rBL
mFR6ClNli3YwfDYFegU57DDFTCi6Kus0gvxKsG/KnzO5fiA9DFX0RsDAxic56HP27nB24eF17vC/
N5lpgBTi8S5gSnnfVMawrziVLWEp1Hx2I+4qKDvzB2fa5I37/GJ75KSkIFedbO+7XLN0ZiQREgfL
eQPs6xJxn0+xXr4hubj4+lVANpFkBemt0LdEnwEI1A5QsCQIq9yTzJOl6aOBtDcRSS2EXAjdCS7I
NiPWlBp9Sx6rdbyVFOT1X3oRGuqAZtYl0eeUiSE1CKvA2EAXWtFjPfNhP0u1IAmG0UiI9shQoFoz
DrDkwjZVI9j20Va3GVQwf73SvoVddz3f96qYdEr0OW1gqUmPUKHNR3dKYQlYZMUDpv6bSFEqd738
35RUQkOpCH8HEyVeAo6tFshoJPR5bJrrz0x5AaqUU1fhBBMBblz8kMFUY+lX2y8KGhVN0sX8VAR4
Hs6fKAO16jSOdY2EdOTKsDaUp3zYrkDO7H5oZv/pid/eK0vSBNvr+/IK2C6mm1rAfsMIpVatF3uS
Ga6ahrUSUArauvp46jlMW8Pd36sXhmeXPayHvozkrGc/AgY1iS8xg7uWLWpaY4+xDN9FT5zpqT5r
aGgWT1L3Kj/hAbPAPkPk2/StnBBs+APqQmJaQP9q+7ivDSrXtkSrVy/SE0XwC0JezkxOxDkD3HqF
rRgD0qAhXPi0VDpatbtSOEeuMBltZJ72ek0A3ZrqhBKKQcS6B1OAMeuhW7Ry+PKfa1CPN998kD1x
TQeEYE9vgSDeEP3DLaz9CAxCEqypVXLtWAY0EU5wYNZ5M7FqEacRjwmyJzWAlolI3bTFLIw2BGAs
wMmAxkqoe1LEwOKbiUSPKYgvAcEyPYG7cQwp3E13E68f+4G8pBNIHHpasOL+Su5OQDcWZT5xTQCL
lYECNL8cvTx68WQiVhtZQOYwsnwaa7PoUSqjueFCVSbMPgnfV85jP/3whzT8eQw7IOGYvIs5yfET
Yo8X136J0APepp4J6hYSWFcWyqCbPcWNOUwqN38TAKfNmpE7333mfy9vttAwcN19sVTVB6rQITpA
FNlZAbHr9Lk+4msy247lX6qU4C6yukdZIeedtReAacxND0kOjJH8j08+OX/8QEXwsdVeUE+8Leky
KLHoLE1GZG6jF0yNGvxU6L8jpf04V3yzTYi49RupNKA65OmsOfDN+oLabYjwjUdTL3GAGGmYgHKS
F2FwUmOVo+JFzIMtyXkmpmLPGZF+p30GjkszU5Dvc6G2T9fulWXB1H/PAFN3RUCAfDawZMPFKSQm
4XuUsHh3HiklJ9Qb+TRRxvsqENr7L4NKKTHARtJL7LlCq/4ek/kvIVBrddRAPQ993p3aZNSPfbGZ
KBdR7Mnhz4LUazLY6OixADYSyY4P4lE5p9avqi7DheTYQUZc62ALkdB6u/gRf3dTbG1IZDl05/Vl
ILYZfUGCzNjnW4C57wh6o0o7C43UpUJJAMvp7qmtF7nK5Il0SspAO9vGNL3vT5fXA3JVNMKl9r76
biQ9sd4WW4dA7OaZI4sZxBCRdn4mAEHUVjggvdpaUmTsAMa4J5WrqaeiwHwtCeb/DyoSoRaicnDH
8bUJsWIUkAfAaNoCHf5QS3Y1TbABD4IXfv2OW7hW+zeovWswtD6u+7I8cptCZyEAau9g3osP5+K2
oi4eyA+jvs0wz6jejxgzbzCxMSdgNrt9+OIUZ26a6RW90DoG+1Yd/HnTQmIwsfB1Dg2dqRb3se6Z
aAxpFKjkU7LrZGs/OvpKNgdnhTRM0tB2jMRR+2N9xCuBVNXFoal0eIkDdrY0XJ4QzU+tV5/7Amal
IJYP1AImuPJkNI3+MsnAUD3WuFcLcKuJkDPbj2xFNRN3yjnPdfUu0AxdrQwesL45hcJTo1oCa3vD
P0jny0tpVMhmRs9DWEepeGV0fRe8A23Ormu8S9LRdmsWIdurMtuZpVyKuVMkHQpWbpsX7l5t/AAL
uwIHSEoCg4MOR5/bw5VFanqKyfSNI8oAJlbHBQUnCy7+nFQ2uUky9EuUOpAC6y2qv5iM+3gE/XA4
GWExCMP4YnP1cf//Boy69S3dv4QfV0Q8Wv4Vy3oUPd1RobOBjNqxF/PIcVGLfIlw68HL5W2Pvder
FlsyxCX6tyAOp/m1nmml8QOWcv5Ef39Wjm2LG4ar+PMf8X20IqBAoDAL4bFwVwJR9qm0B9Tv6ak5
4fDe2bibxJ7QGjN6L9t2CBz1p4P3BK8OHdTZY5Iw+2QLiIYnVIg8mjeT8PUiCo4N/6ejb9z5kGh7
0FZ0dT1us2hTPbtp3qMKjI4BXaD3I7SugvJgibDmx+AfmfZWWAR9S0eLmcN1n9jmUWVMSlb/Nx6k
S8Ij+nS30PLAZaRRLt3oHfL/DjEH3dzMl5/dLpoy2F+pHlEv7rDsTTPgM+L0N+qjfdx+SHoZ69Zf
VVdGKofw/Jy8b2wuExVnr1c4paykoDFUhh9iXp8RJhqoWfkOjmO9PUyq3w1XDnSL6PWcDzySUPi2
D0gjJWRhw6hINAp+RNQ9+I9JgXDLrfuP6/tUcX+nfrGYFYfmfz0Oplonmzpi4WvSk0LyTQGBGI29
3QTyu/QSdbdg2qeGMfGm+WXDWBpPK1XrSePONNW3qAxdqqgLLlFELsyMvdZfGbSgG2kjNjGxVNsK
w6rry7bD0Tx/f3xiyj5lihyZODwwFfKSeobxq/UsS8ssyf+Q1l61ms2yptYMEN459lNV7dKfAiau
1w02dL9YiIgGaD1PggNcX6eSr8NlMnNIxbvUx5c6vcuduA/JX/zOyNAMeaIxPNEjSWS1ercPJ5B8
DZOecE5nNplNXiFlpVDR4sSIWb+Z9vFHXsC5YRXSX3VcipMCNsmzYQT5fhTaDg+x+tsz8EX0QgbD
VnGo6gpnMiL2tCA/hU59UgbYdrltoPRFF5P6s+0v3CRJtexY0m0h97iClKmeUcr8sUjSZR7kktZt
mbYOG0ldy8C0WJ9NKP7QFpULlIrOEHwnAIU3prPnaAbdYJGY5aasbcxEoCJ3GHHZ/tIxGyUuDwZL
GqC/FkBhVUSae/vwJrrhZPWN/ADFYCLGkIi43iRk7jrtEFCICHX8QVfnC7/T5kbAEJJf2vqBIF6s
a6spRb5uuHAELqTZ4I0ZJJl4jhVCamPCfWu2me3f1qdtMDuvhX1zCm1lCm2c50ABdTCa1TqY3x7d
LvvGy+2wE4SkrkHV7nMFNQICeUFlj20j+z0UdzseRoGnX0WdOa1giJ54ZdnK374bFyjOnqG5uTyI
pUiuzA6xBCeNtj0ug5izaS2R49V4SG7qAE7Cq/+moOTpT8OR3parqWk8+prRbD9ucJQfXpFWsSGF
zW2c757o1HEb3ws7jRVIe/g+aCBOqp2P1nTrN25oMtuBaB077bEdy4zvFp+DEUUb7WVt28KwKpxq
r8c2lcF+CfdIXDRBuH/At2LWoR+quBkPkQogVwPszfMfnHnjy5UYuUZA6YFFMISCnAFa5tivhQ6l
GScs/lEJT3hUSiQ2GkGUR0hgU3bkqpcxHlOtcLkgTK8wahUcFffUBTS23PUn0lhdNXbzIirXcnB8
qM9RhWvbvVa/KzvK68OrZTzfzmtZTIUqcVt0IgAA7OtwDIi8ihkaUSklpkEhCnM+SB8H0+bDoyV+
lTRWEfJGKK10YbBoY+CGwzJQaXV8S4yvRTNs1xTcDvtHmxvRAhyQGSbaAw/8GWrcnBKvi6P4yogM
XssDyBbge1SYXs+uWYAPwfAButrCelz5kknKfq1SF1WvS5gyq0K3k2AII1Do+hKLeL0tsr/abmhC
WhgLiI2Lc/BavHphT3rTw30x6x2L+TEnv0df8QttvWf/Xn2y0Tk7gjzrV4l9HSbJhoMt8AJa8X/l
ub6eQC3upgRMcwhHhjyz9BMqhfq4z50UxvK/FlqI3O5DcSB9V4/VpaKpYbnLHTasn10kZFMKYSPj
shgcAjiMRur523c7YBLheZB6IuQWGusgzY8G/4tNXspmpWmgKKtQNkaKjc7/Y6FjlZ2B0Ft03O2u
uJeLcyNvcNYpD3OUqwm1Hu2RyHnSzd3CC0PxNOhvQDx9vsBcsBZ7UjxY5hi1YkaQu7NwafZrpQ4J
ZEvl7UAKv+DXo/9HS5F3lRmWP6qBftCHrgFC74Xzk9XWSup3GpMENzAtBaQ9yeWPQvSb2NSJxUVo
BC/Mm1Ic0l9rSQowfgTw5R4s09xFzWB2JHSjzNIcVLLe6ElauhnzGvze4fipIQsdnSYom2kNPWkI
iI64MyXT52kehxhIrVzWPeryVkiLm4vWS/B639t46hPeZNX2BGykkxPwEvPyqT7Y7pfA7rZbxK+B
q54JZiJ7MzHR4lpYLRc/w+yfniMGZahf2ZO8cRH074nn2QTL/25nn4tlugj6I8w9RwYxlB82gajO
6eOQj++wNUaS5Jo3DTfKnKOSFkyzzqSNV/8j0JtsjIsbqcsjFK6U9NQ9DFJIb+3seB+ekmP58xuJ
iAZ24/o5zpK8J7lv7W7FaMnC7xOyMQ90XthAcFv6LukdecCY7ZCesLGhkwsz9owBAgbFF9buLR0N
w2ilSeG4lYCfygxtdjFNb6j1Du3xWLOaAaGxOVVgAoTHyhIB+R8lPuKgGNd09a1baqwiWNbhJOGk
ICiVeBQOD4uwvkhGr91kETMzRYJxIHaVSrlAOI4JfxJG8Dr/Vle0Qo0+cJWvcLJxoCrwPHurAExc
IC0HwIP1XfjI6jOum3VPxeWev1qZdRfQITX73nq+5PLtTtoeBHWDqctft9rOKxTPPOkOwuEXndK7
0MaYsVkkLrYYYz/0ItXTn6SBS4idIxruI/kOQ8DH7hJPYThvVEzYOsOPDNOtrf6SWYW5viVu40fm
1Q6jChO3GfX1oBgN+//k7pWLpxKa4yqKcy0+m1FoW8Ff1CSMeuZ7L9Rp9NHzsNZYUyx10FCrHBaF
yNr2dWO1LyG15EGKaowbdWNjmIc5mpNsr54C98qtzTXVo5tddrDGnwNRMjLhd29r1/w8n3vUvdDe
cY9s2n+RT8y3copcU9FRLJrJ1Y2w5bMYFZt35tEd6wPJeDYFIHfmWdiQqgbgrKsnVnhPZlp5dOgj
OFH00Arlr6Pb9XUwrpYxJIQYI4myatbIxIMRq4DtNEFgvf5q4JXKksU59liFW5T9y3Px9Ki8fFFP
CpNrnfPz4WrclJCc9yl59znU6YynHe/MYytfs9gD01C4z2ho68uDlP7hbAW3+AcOcGLfTP19DUii
nMzQduJ+ZXIdDnAUW8qegcI61EkRd+jnRpPcbhjsbt7De3Kkad149hqJjkIKt/YITZ6d73MM8Arr
nMyFDIp42+1U6R8EZwykNRlF29pGJq9zQ1ZYFxntbNRccH9GweujAUjLX2m49oux7hSLwbH2vsIc
zncgeVt9iZHMFyHmGCPtaaVMovRMDrI5bUO0E+nGh+ZuWxt4a/FHmLwY2fAQ3RcGT/wcItDUKXus
ElbbYYb6oqKrQs1y95WLApuMSZ5tQpDYMm0F/btVa4qIfxg2d0ay58ahr6QZa/FUHCcrIXnTsgl/
DxDjjELfke0VOkzb1rVat79S+njRthgJXMh+CnpxuHSxnJe9yWXa8NPURFzwRpzmrNo3wh1S85JJ
mm5sAXKsMCDdKedSjHXT7pJ9KEalrzgCkGiSJisIKQLO5ltf5I4TDQPhyF/YABXjTmyddQyrVrh2
0y8qnRZEHUXYN+Dw2mmBBXK3VO989WBasuNjvAdBTa6fNpuGRlSmW4hcmiJ5IVAa02sOPJo5bnGO
4WV3ppSQ1ObryD91lcDNR1mTE4u3uwbyh4oJmicpcIs9DoMmVSTNoNiMgrh4NXbXiQ4dY30Rs7m8
izOHXeClya5cN6ic6tL728V4EyJx8jUNL3BOkeiBdAiNPbZi3IfwlOiAlDVNSJaFUU+7u/Tvyh86
PDMsaA9Rs9VsJORYHM6/kYzk2bOxCLfoNrihQdf0EXSXqUyYkZVZFiI/rOUPYyUPxdR0fuIJhiit
MKvDgxKDDL4XfDy7sS8JLhfgJ+1vbMMW33nK3fzVPbAR6LIen6JxL/MkISN0Rs/v4b0L3JFVhmXk
/OlH1hDyh+1J9zwjeIW/MCfxpSCkW8z8AAoNO9wA1+FChnjPrWxvum90jjBU3SCDD/Wwoqj1ya4N
YQuJqKjgRy72tBvli718/XerUnCnyO1pnKI5b6v0COZP5UcsK0J3la7okoy4tkcChdfyq+h0ZqcA
3rCc2fbB9SQ9Pj1KGh5xr0YWZXwVP0kTUQkGXoLYq2h8XLiDDy3zOmjSS2tpJd58ZZyhsXOPC4Q1
GQoc4byf+mCEuRKtME6ZH5dPI2h9KGv/KUqXYEBR4N4zHFptlD7TfvSx2hybmjHsPwqGgdvgCUEZ
lcs4WqEgWvXZV7SS5w+oRUTNX7vuOnTl5/JJEaByWuq54W5IyWjbX+mHchXLkfbkcgrAP7CknVuv
f1jZb62N+ZKfkYf5WnZVE7G34X2PT7ch8ciAHi84e7UAcKdZXhPCI/KxSNob2wtBe8huWn1fQgHc
KyRTS8qSejPl2ILRtsNL0Ow0XSKYrlWJmIyXHVOZOA4WeuffLelYwmIY79slAiGzoKphMa6/wYui
mQAIyoLzFdP0vozjGZuyeXCSA2BjRs8frmISvZ6gNeQP7lvL9+nkSMakzXEaxAldBjHShl6cbKV3
QlB/T34haClp6NrxsB6s3r4tWDeHy03oid+WAtmv7/Cu0n9ul6YLquFSY9GYgQnApzi8Ngwh82d2
Z4eWJkiXrBpUrHmDat9cm6ZsMDkDhp3Tciaxd/geekPVl90fPP4/3LzZ90nm8AQFEpXq0f/UhaoJ
Hc5rMyU4O+0tHf4LHgoptXnx4eAOuHUa7NsHn+VvbIO1CNPLFODgH/IVrDc+zRIRm/Ca3DUDd6hx
6bEv0O7jZUBN3S4+9e/ndJDidMqDNo2FLVuOCJbUlpojwFjAGq4Fj1tG+YOsbzi8ek/QsSx49k/s
VgmLXKZ4xGezSL5GQpaoVLv5ztZUkTeBzY+ANTlO5EQEaVcvlbUyf+19a/jFwnKjADy64i+oZXBl
k5f1yojgACQd7vM8P9hu4iCIGq1wy5lMb3XuP/g1swPDnPOpuoQVfjGPRck0lXHNQ24m2zbq5ZSr
5/mOc+nRzCPvUsFQfWnIqXPAtiT/awlufJF5ZxwNAcrK1CD+nUuJdnIWEEmsswy7oa51FjXeEmB6
mswyrJWM/lzmFK8RpURQ24P6cvvKSSnsubuiy15Q3r+qgXoEoVp1Q8i8pyQ3m1c86dP72Ocafrtz
xQy198kSAEumnt8ZoeS3gcMIYeZQasP8RrZi2YAjS4AOFflR0fkG5yPrGNha1B4ZATYtbc1wXUnz
pHpmHNsuiDTEVsRNuVlqLpIomTkg7x88f/cxAaVFWbv0zs/AyABULDLeb72awbSaPoA5dcxtiIG4
fXL1WB3p4FrGbU/zLYobwdZR889mxCW2sXS00lE6hGrHGzctYCZOWH5laAMtqAD/8ukcrRiDy4OR
hN5EM3xRsOlGEhHHtbwoxyKkd+zZxjPzncNniA63kRtHI/qbywT810GPvf/JWF5CtxMy8/zDXdX9
j1zrpJCcLxP5KY7/GHLOthH5kGlMi6n2mbaoKzEixwkzQz+igIbFTvsiwiGvN1acS7Dp7f/6fgK2
iJwP0rMP0jfKFhKiqyy3RlYjMsGXqSvNPxqJgxvLk1tJbKj6Ho5aH2UOZ6Pq1+voh+zZ4DF3nbH4
4Ih9qSgpQMunlkyBnav8jsaoclS+btw8krZFwFNsmPsC8UKf/qkqicJzLyWnqyJGLe5ewSzNyRhd
7VhjBTo9EWTtpnmKtHgpVCHwnvo2JMSce5F7sHuPyvFtCQCH8lBpKsq88lUG+t0QQanygpdcNQj6
tu6nILOBo09SjuyUjWiG6moF7kVVDx5VOne7fW91NORro3ZUxgVangIlzC+g9n2Z0mEEsQIPPsMY
dWe/xxVkV/MzywHZu5ioY8ibLJnToae9xmDB2M6eVwkJPlFVPjTxnOWthkOrRU0X7KA4+fn5nbj8
Up38QyEEk0cphlbW7RLJm6jR2UpKDOgAC2p2o5JA3W2Ok6fMFfVcYywhtxvdVp8oUj7DHgFdnMFE
aRIePVj+qnQ7UgyC+gTXVjd703dfRv9AIAVmoh8jWfanmG5ssxP74Q+1VNegZ+GWfkhjoEVB/0yY
qN9G3qJrLBSPGweh9eE5LHEpEeLPD2GJ8EtBQbEv8DiLEDuzEb04CaHSq0zRCvChhDEWNVeU5LjE
pqOyFNjkXlgrINqYOUzn97vDig+9/u3bwPhDyZ4xVqvmcLa1V3HQtqf8hfqJEMRK52ZtLWnTv4Aa
OEys+Km9i/lUaY+08LC3fNJ9bXoQpGRBhILSfya2ALPHnxtAojkMni1zhfT9W2IfPXu1+JfLoaAu
uvUR3EoHgDgQA2yBh6jHbwPRcS5edf7ptrJQsNIk19joKj6jSuBmJNKVnc0UqNEaeBQQrNnJRA0Y
7QoRsiTMyoiUH/cnuXakeI4NagdewnrcT2u7O9kRdMfOUhIVlsSodFvZaNNEByrw9+BB1bddSEBJ
vAStM9qX+cPAsX0E7PAJMkJiUnt7AkIcShPcnCnub1Nrd+35IxQggUyDX8g/JdpBxIfUQnwwRiYA
DzWUgqsDoKz8dcPY8aQ7RDBpuS8zJwyjnOTkB8mB4mv6VY9m1vpHC4Lb5vgLT73tS4UJAsiDS0AH
pGjdnDvA0kJbeD16P971tw3JtHJaIT/MO/gUB43nSoy/jBtcFkXRPZZlSmDTQzXnJNtqWPdkRKdG
F2xzsNRvh3C4YnrD4D1pcJzQNESZNI/a9CD1EnPPZY8TtdCKH6P6stEpESJ+ReVyQtkLw2kKa6ai
gx4YxdfiXVLqD0zAuo8pKjRbU1ZclFpniHkArlSgNfZihgl+4MijEgHcIq5rsQ5c4h2pLWyowbUH
c/kMMPFm0fBMoiPEuhOIRk+dncnvecBqfRkWYi/U6y9JYgDrzzIJEsSh9L8hcZ3opHoVLJRk00Zu
PjgqZ2LKpQFNpnUPi6CqlVNNtzrfPcz9DENFrncgsT0pXKjmrPKGzZEJSJI1C7LIrFDcys7Yonjt
9u2PuCgCtZYNiVRnMHIbFmxqDhGNs+tgpRxQWRm/AZjwjZGCFc2dBalsKP4sq8e6/jpFbrgGXWd+
GBmptfKxfIfERej+zscxqqMC/j8LvS6nPU+VcB6NpyNF6GtOzNXTa5xSQd9yo7V5eq+4hecCVPBV
EssWotSgkauDTQD9oypVev/MQi66rl+iDIwQB6VNBZ/uy+l/8C8RiNqMQYNBPhfNVmFyqvvv/N7m
NCfo86Y/YfN8AG3dBZ0tlbjhWxxETG61tgso5ozbDo1XxzfO++HV1WpZPz2UnWZOqOCkGDfkA9Oh
UmyDvA8xvyAvuzJJVG50MTbYVgWFiLUiwK3G4S3IcLKnDV0r/GsF7z9huST0axuNBxzRsR1HXc5p
omdY76j9kyZqYtrPf0MtzeqwM8UxjjvlW9e0AHkpgKbqIx/CqWUR5NHhhN9I070w9sGO/j0fJgXK
j3lM8fj3WXe/KbON9G9LnpfhaOmISW99RA6ewfvr10rLwGg8NHM0BaJEnCHWq0Cg/DAH9yK4zESt
Y9R+YACUBmryoyKo8VE7PkMsw8nZvB+6gBqENbxaIyTPYYxBUwaUPr2E3SmxRSX54/Q+XD0XqyEE
0rI30meFmniLatIbLXvHQPRj512qW9JnT1Q3arzaOGzKKA3XrIhDaw5QrOKO2pAuSkmQJaIRDF6j
NOuwzuE6saS6bOHU2lLEeqtkmVc31pk15Ze6J1RHc1pAlHoevl3Jymw/yGl0K2YAEi0lPBqVWcJe
pQVh6UTL4M032nni3YIHGhu1t7BwjUkZ7pw0L3opCma83Td7U5u2YtUyRkTXDhgPTJlL37KtKP3r
KHDTWyrFX15XQ7peU2QjZDCLlrkyodHS89HgUTcxSJELyr/I3pdzgpNc2Zvyynw1MFgdddXmJOdj
VrPGtwrrnf5enH3UGxenspOak/aP8xmvWts2WWYMgN33/UC75izy+HVg0n+OHqJGb8EF+35MYTeA
P8LRIDzHNfirPNEIVO/uOG1yJ1zlzpDeGqz7UGXnjk1WSNIhYho/zMa4HFLB0MlerazfaEuIR7Jt
SYpN5neHXoXA6zEnAJU/NQsSTjRxeanANVDxzH2L4LWgaqNgHVh9lABBnXnpkWvW3kYh+7bUUNwH
GkSmf+EOhqiWIIMPJCwwtqjPpY2CJGFLyX9m6AAkiBXsD1ofEBiHrBuuZJKg1ZY+NpSWT6fP6Gm0
RP44Nh+YrMmKAh2464XlJJPQx4HhqssXPWGh3bxrB6GOqdRdzGRT7D0QvefHdmCC7uOq5JgNzJoL
svsdeOfaWrB7N1SKBFn2z6g42XLSBo0AOMeXij+ymAThBNu1dQtlCvQvqKtD2DaFruAlV8Ggey9o
Wty9loXThZdmKpbQnlifrPNp8UGSd1q5Av8Pjw1ArX3dvIaH9nZTJTziVmiw5WYQl8IJGZ75Kskw
036VZMroA38jSzKrHJadWFS0ce7tL+6vVrlLg8SECzg6NvHLf1rv8v/Wuoq1hEj4Mgkca8P2wIxx
FdZt/RRuHwsrqeUQyflwopOIdidhp+FsZgQG4NNFukSw1ZrLk+FmTZhGDkiz8lXtX6V+IPJkjzau
AvImlvEUc+bpy47sG85N2PAjIYhZnpR5OUK4MgB/P/Nu5mrn4qBAEJb+wocyJstfObqCKTbFczmM
Hb/ml6bCMGEq9eys1RfyXtudoTO1iOfKFcpbrlCBJbFLzmt/lLx5MLztm+8rjDQngBM6TbO0nsFR
i7+dIqjEzGjulzUQjEaES79oZ2V0NYm+n8iw8C5p07kEJTlyioSQPHXVVDmD8ICaxr6N1FzU3Gy6
MO/cNHmtqAuHEun7aAeR2VyK7aT3jXMGEpjy6zA/xZG2JjMxQElaIeglpvb/zrL4YJ+IVFKGKWcf
SSaQSurfl3JummNZN6zRW75f5oxrcO5et8YTIxpTmLn0PuzRXbwkx+cpYC/6ITrvHcZfseZbhGRj
Tmt7xNoFJrH5m3i+yQexXMjEroOtAOP2iYVa8HlkuRecrdh9CJqX0GmJEGnZ5AmdMOYUz/aFbQtR
ybNG3ES6kMpJAvTC4EAaKC7HrbCJLNkoN7dn7d4+1nkHrnCMaA+3l3vQdJJVa4cBXvV8IHhfZwrq
JAhH/DQeQGZmI7AqD7w7lzKBJDSKKFsfb4jA0QUgD8CBrm43SR8yleKpw+lCqH45CpGbGWyuzYgY
PMTgH1AlxE0pNPsmLNbvYb3xLvsH9IAfO5TXPGu7rvkMaQoHqxM6Bkl+yz8IhNgXXXwFnJn8wJUw
ngNZu+Qtb7m9wuo9ZN7tbfrSUTarA/06UBpf2HL1vkr3je6miw/B3NaBo9xknVFFDg0QDDSWdPmi
U/TA9ck8iD9ChQuxgUiiG4BV5raMWPm50PtRXKqc0IQw76Q/GwuSa/+Ch1tfdbXUJKezjQrtiTI1
StZkhp7XJtinDMqbdkDVM8EQkz1m15Tk8GqlyM79Z3IwEPMzx+otuyPBXfiIl9iGQDX14PzEkm8n
8igRRSfoZeyScIYu2y63B1lnNd9+JmFFGYXm0u7+NM4x5TU+T2mSE1aNtjVVfq2QAcGxcFvXilgU
ZABukyPg7MkdotIgbmOFJpl05Q61iKUTx/g1QMhWNGEkwnWkkD78ihupGfXTSJlOp7fjUU0QHloH
8nCTR/t008iMaDfU7Gs2yBH/+r23ATEserrqjziNeXlrbWBOvvB/aS8rGar+w/hfQMh0FeM7xEjE
xm73nn8qWAVt9jBWlnK8tm5YgpED4aAUaRCAUAtc3OOIBW41gJPimR9jh2qVhhqWJjDC9EUImRL2
asaqPtBszXfOu/agDhZQJatU8sWC6KdKhnR7en+tVG/g9wVw8Swgh4Qn2MRt4cs4cWXSHNN+pS2p
8MabHfmvfvzeDjh26/TzGrRd7jgl5pWrBz2OVMz8MVnvm2xQ2soL99FmY48lQfcVSN4QSf1Ig14T
ntqD6c3aieA2yjBWNR5H3JuYa68HLkw0bEw8aPwaKIMzN97916NOuFt/+diM4WPeOxxBK5ga71WV
bMreZbFBkFQ889mzECNNG3JIRz+Ui6YWKkWy2Bx6MINki9nvZOe27yf9JP7pL1aqeFy38fIlRVmE
w/xQVQKbEZzAA962MzFBDfToADX/Vnu+GBbxlZcml4XKnVT1k1dD5/aIrEzd3iNjB8J6ELqFDPkc
HeONSnuO1P+CVf3ZXFbglb6uCMdtMO85d9E02B3nXbQLUbj9NNeociO80KtBIN9D1Pph6wsTbIus
qkRYYwUoPduXqEZssdSSo3XP5lzg/o5HKWoxnZ2ZeaLAjmBYi+s8yr5Af2ecR4WXZT/dLZ9X7y16
E723Zemwfbp2ELJuyVf6pl84l7e1hnvntx6hhuZSNWbB4N3ZjY2jpemzqftwivnSYzRxe/wNSxt0
3Ecex3Dwxq4pyYGvYsfvvaM6iOQBUPYcTCHdTmJv9KrOZXeiK4OTPsTmM0hgOUOZSL5iyWa/hWaF
Ln4nF1FDDFBnEoHBnWbcvyyYsGs2g+vYqT/78YRCtKhlsC3oSco/wTZQ7rmyZ9n9/Yv62wAXcZo6
kAhm37TR+8qONyBik9zjnuNPSA/Fr7ONgEPAn7maYzMQamZ10TY378nkBDrufszQHpjipw6G5OA7
0xSuh/W86k0Rn0FjXCoZYBFFTMaKZiWEYBOP9KhQ7uOGTRaL4VNuixA/w2H8LMVdaqje8g6GOACv
XBU8E72/sLJzxqpNheK/dWezoI8iL2FH7tk1FTNYE0q6l7Zo5dpD/CsJ6TMxbNuo9JKS5P9Xwt0u
tMUJ586wTFg8TyFjcVg+jt+TokZS6bURU4OY2YX7/LnzgqGFQ6GCvmCkcyyA9U/sGiUQm34wYOvl
SCysYzTSnMx8Z3jKV4URdJOAoCAu8QLWGNQPMRPTg5Hobp/pi6BLWWDbiGQVWMHDevdz2ddw5tFo
/3AfIlc7Fwon4imhvqTTvm+DQ6p425hIqrHUo1n6bdT93BjDDI5mD7EFjV+QrsoLO4eL4lSjuJZf
fmUKROtcFPWaxeVMrCwNjviEwD44V8nJnEsF92oUPq1HqfJP3CULL8ONVUSpuBLBppKEOohfv8sT
jBi/VpHudxtUkQUq2L2qFtdEroKnjh1L0Odk2nQ+oaDpAKq/Iw6xRCihEvIFnDYGoogtP1dBTyUo
wgdzK2ir6XfqRw35KUVXLtGrlA23+ioHoDtOlZ8Q9tWyHsy8wk5yJKI8JvW+5p3E1Ij6Hwg8nTL1
26JMgdLpSqHqsGVKtcbN6va5CRckC4UDwcNMQx214LAHPOH5foXgfC+GpPP6NNfoj3QtWB7ZVRVg
y/Ti4yepj6OfGxHh1gqzHguYz3bVtT3TJnOOitBZGOUGco7bV3L7DUWwg5eD5PEIQqN8QyALDRtN
S7sM6P2Vh9BgvyT2Z8KB2ZQjOv9OEc4uI905tAnvqbVtS4J27jps3J40Fyoq8kQZm1rUR7Ig0fWL
XfP7Hzo/uUUwyGRhJWiuWWl4itkJq2Ak5P44QcJ1RaNc6v9/PXK63+6h3pjbqRL7+ww6dFJBRcU1
sWexIR1+eaep6RSuIt4pBpN51/afzgRV8qqY7Ah7ZQN9/SfltEaWO+0muYq/i+0jUAK8fb03Z3FW
oIsya8xPWtuQ8hquWLAbUXe87Hq88T+kqql0zPjRSYhqQokddigxbRZJR4C30y2xSgudZmj194yo
mop8knSEgZ6SYeSufzX3MDvZPuC5fhNEbukuM/PtaetcISfj6UluHTGq7/1MKLVWJGS2Y6M0CDWV
KccRRsV5hGa6C/CBmyV3HhL3uRnoTIn2q0EicjcP4S8YzpxHydrKe2EB0dRE0Usx+inUPSoJ/H30
sZA7eJh9zNrlcUxkmyuf0+i6qXuzitV2rQgUG40cGR6wLHJzebmz6M5dpojsTvswRmjxEskq/FoZ
dmEhPOMXCJHTsGOxmEgqF4ItO2LscMGslyrwTuB9y6gy8ywrfcH9a+3EzHSR9nl3nahiq74J5OOf
fc8PgVSljsEk4TKBpgStSDDFEjb7dG4v6eWPfSqjRCMorwTbcSvJEuNpiz0qttUlsbDZrARrasC1
K91ZG4EYwEc+DAlHk0LJLPc3gLrDxewJIg562BfMK7WMmht9QlxozpZdRUKGDHIKDNJ0VscP08YW
4Hno1Kbl6GbjdLKDtuvYwcSJgo6WCKKSmR/QqKsuVojzAUKBuOH2lOgBNEz+L51MEQebLaCU7UlU
YhdLUtMR6yu2Sg54jdGIsRoqhBlZE9+UPJoKt4GnXHb2H6lXGwnsLeowmn1Et0rO1Yqfu9J4EObk
w3W+hOIk/8fGZIO+eNsZDvvGfGuUZkp0hR1WZ27tMMASmx9t8nA6RSiR298Q2L8jp5q53q+GF2/y
q2Wz49984Tkmr0Idlzc7ldkKqszKgoH0ypMMwSiyFUj9aJnpsf68Bzkbm4gK8x5hJ6e91Xg2MPxL
r6U6yR5Vs90jw4wObQffJPF9Ip4+R00ZVVBs9TPBGeNoA8h7kDX9byyGqLM2z6Ug5JB70eawMgvG
XxJUdGGq1jmlhQfZib/lB/bBV3P6gFwh61PRbXp3zkVrSjC0IwvXO+/e/4L+2sYZD594bDY68uDI
iDpTh6pacl1LsvVB5jkIQ7Fta+2SV/ALNFueRtW1lBmzWy125L61NaXGA1i8rUXaFZx+vKFH/Lsy
bHwJB6UMxCBndSBe3vesoOSyxal2NuvklUtWmJaIa7dc+59qrfkMT45xm9uVV57VHuPexaXNJtCB
34pih+VZaz31/lLPTs1GcLKfux5pWLFUvS51A1LPPVB7t/NxTZunME+G5LiVoG97JlFNsojOtxk9
e2HBR5d7Gr6YufDiv+IQgSMlGgipqhXwo3GSomeWsMMbs7alivSHQFrcowbkxEjU12/vjUzk+zak
bOmeXaSHm0SiHQFELmUh1dnNgGjdsnmL/WcNPA01m4HVIw08s4526cSPYGx9fiGjOQp54882K6QZ
dNdoNX22bbWvVQvEZs+X5eUkZiundev7NbomIQ2ZRkuOaTdtkn06oh55uOps5nkQdjnmEp7C+HZW
lm1QAP464mLI9RjCOz8FtM7OCvuSgaAoyZ6+aFfBlkuSDehfyK9/yF+QgaRNTS+/9w7ZtZCBuex9
9wSKpS7LxYQFA2JpN/4IUwJS9VtR8nL9PTV0pzIjn49y3frtl5qOfViqZLZ6gF5bLDg0ZHAsmP2A
2K/nAwFroJ6wRp5oTHVT/tv5PtVELxu+uPOTfosMc1v0wsgDObf3k1053WU7wjC3D76fHj+fH5O0
hQw9mK2vz83vH1oa3M2rLCwYiklcUt2EjqUWORF5L5oL6AsoK717Z/nV7h00DRkYXdhN7+uUOyZv
G1Fs0pvqTInQNKgaGsJ4q2N06ReN9IBSc+tJ8xNegvUc0TeTGei0RnTH5d5zPjfswsab0T85tXC7
Zsbq600MrlbSBlb42V0Dl76AJjkf8olHfMuTjsnJR+9sTZrTLIw9tkn46ncRjT+k4TEtc0j6pPWj
qUX02oLyvWQDIGYlAs4i2ux5g/2wz9KowkmATFRCNisbBVrPxeIy4eKLLpmGB6kR0nc+O5ywj42A
Cav+Fadqhx6oXBjP6XAkvJoMS7Mb7nXhFSVbRN81d2NAtEtsI5DeqNtgaD1AlzGcQIvShScgFA3d
H42Di3rbbZ8jg33ZU+lH/f5L1e/w6Cw6cWNkgaU8Hgm6f8yByJDOiWfbNky5vqSjx2mXljpLOnwS
7QxKfqQOdMFj67rZVFeQ6iP8z3MpYQVwnjN8chJn6hFupKTq76+u31nQB7DyxA8R1t6ui/Mo5SLb
v/LSra1sjaWEwvBZEHqGF1PE8RqNBlooAKqTMHBAAmVV5+9aip/N6z58E8/hxThvPIE0J1mAVBDF
siy99/0d0r2X1eGIPft3U3aaBS9lhkWNzKD+TdsFl6Fo+tpXs45BTq6pE9pcnpfunwyHuEjP4w7O
a8Y1L5T9GEQc/GV9Dh1jg+zUBuxXzEY51JblTqsq5Lahpxo7adHXj1/wjD1vk3m7rlJD28XxvHlY
8ttehX2HxDquUD9gSxiUYKENZ491ax4Yfx2CqHcClW8Yao4BRA/yeG72ZanQmLnd9nxzDbOzCyMW
lBCFSx/pdBnUfOKAr2rIqCdC6cTetd2mAgxDhNVjmIlA41DZonbc0mH9cN6AM/VdKdtJ850YN6UR
n6UuRpIT6HaOTrP0/ludyxrPxEkAG0pJD0C7ZsOuXlo/lyoMno9yFKChOYgtx0cUsZNqod3h7U8J
y9oN165nVZfpBQDRrzZM/bThMBf/WTyOMlcIcXVPF4rk+MfsFYVryEvWoNZ+6KgUZNCyGK381vbi
wkAelgFc81F12NLTaD6SdJqApuXtgq2stlIgluHHUbV1vcn6vxR1+eTcUyV++7m568WwzMB0rhvR
PwBzENdlcobMxw5u4FPrXKtEk53pa2aC0VAxxZz3Eq/UttNxn3rReMNO1Fq29WO0K0oO+ilqQMxc
K7t7jQYzFtXRbIwcxR8evhGKQs9FtHjZDnKC1rtfjvqtM5KT4Qj8A5rfddit2/tVvJhZJG/1nEuC
kVUSuyqBEU/c+q5rNlM2M6jUyKgP/S5hT6dWyJxTzsK3aa3VG6Wwem5DsRpf7UE+j28v04LuICxG
Td9vTNKgni/10/jSMoxqWkV0YCncNYFSt1E/49AKENL4+8VYOAUCLd4tbu+ZhjHbMN11FRuQEERz
2K2W4NOTeS5JB5zVOg+YWYzNT4/ZnDDhBJBmAJEajDdU2raXHj/Ll1Zn27DgD6wCpTBCH/y3cWn3
ClUllWwJ8AVQ60ELQqJxwH9jcr0mFgWHEMk1A69xJ00EZ3sGcmoPX+sHGT+pxfxFhKbHx39bEzVs
UIXHQlgoGsbIuMnix5fTR7bDAzsqlMJsaaD3pjOeEAkS/1bmuDE2DxGSETqLi4V63juGP5wDVAkX
u+mNVVm7qnck90BZQK+qk4wFW0Gvdh2uoiz1DPxy9xk/xRLX9cr2DUIfO5OyEdKyj2SGmZnicNbZ
wG7wKq8uVRQYlCQTtw9fjHmy6uPeGuWdaMhONLgSTzPZYf3YW6NUY3htOvsLIRTdYE6IuzaxKslD
vI1r27K9DbUxdwWOBRrSDCWdxAqt2XFNVWPI9Qsv64xNGpnfWt/g9XFkqIyOw1N9H2629oF/Mki+
iVqQ0iq51bVIesy1Tq7bGddevx/RB5d4zMSA/1sR/Vm1rVH6PnA+4HMMRU01ZGbCqSMR5acVhiB8
UzTeG5dLhm8BNJZ6ZkQ96fu2cXD6pTZxvKaO0wiEYbkyDFcfBeNNmOl241hUzIl00EomjNJUEoct
1ev+/6ZTZrzenphdqRQo5YYIfphKKrUmemBDNP/YwfI4sc3SuLC4lT0kbqH4PIK2WrxIiPA+MRay
+KcKWI3efdY5LnCjYlA845u/QWaxw5NJki8U4YrILMLUscUZfjEjnhdOaIkFTeM2f8JQLu+Qfrch
7AdBl5ERIgR9CBp1ip/kCOv5kXuWw1RhQDxt2usyaHm2RTRvKdLSZh4l9DCjSqXC5LaixsNbIQvs
eOUit/vy63Pav+56iYa2dNtZGL6u5mpwVdvr/u13KWOClUJMTfqE2E4U+AaIcNr7cxfMkWDxe266
FEqzpMRgLCKgDaeky02TnKb2Jx75OYJ3u1MwlIPREv9cjqjMhrFskK1a7Y6aCSuH8r3AdhbOtLf1
6nnL6PxPJYm6IbwhKk/1P556gx9Hlx+3Jm2gfAoVPcX0khtMKNTuC3k6umlop0OtY9FjNO7T+/cX
pLlak70pT5GX9KvQNJvDGATyzH2JEKnPv7H8jQJmDSfkD3FU+q+QmhzcnzJKB8CSagmTO8n0Q5ex
SH0kdMI7oiEQHMZhKVHT3n1A7DK40cutmj+3FY3r6TGZ+GkpvyFigCEOxXWuJYI3wfpnlb4NEPMR
1nE3f8ACNMrU7Wj6e9xuozEp6eI/ouwAIJFB7kVCUcw5GXneb4Ans2nWbR84AkYCsvHsO/6VdEKC
53qjI+dimMvxtA4iEG0GRbyRGjC001Y6kzU71I94MrbwLNJI1QcKt5dmqlnbRVpjv8wTh0DFE/y8
JMWpkmnNjAMMsWDjCe67bfcuN4RXqyMfZoLqHgMGtYdNSBYLEV6QQRSwa+hmrFMwO4vYK6yR/LVk
h2jaWSNzVwpqsS7T4AfPM9NQSDeUwxEYfe6KHMWDq2wZhZx8n1qcFv/O8UK1xe9TLsackyAt/WDb
uBDuLC8ooraba0b2Vaby/v7yqVEGSB37Clxhog510ZyyCDSSjma0d1MXpJzlszVX5tpnh/J8Zd9b
t9oIQtAxPrre5np1OBcqQqRyiBL2cc/3aI3de+AKqb/on+ZsDitURjHPQJzp7cpxvizq29L1CBsq
gkyfv3wAFd7EdjMAJT7bkHxD0sQyysNdHGkcj6RzrNVh1TWRkP/NYE1EvUCuZ1KGR3dwlUj2FJy8
clXTR3XG2gcaEG8/waDLCnN9zZ+WGf9fjwqj0bSO7HimpkjdWFLbK1Wbwx7LxXIdelmHcgXExR6C
1/YsREt1rNbKf/cHqxhRA/kI+pc+yLL74DoklpzeOac8E5M3odnWgHU1co+16COp6xyr1GxqJYQi
iDLQXYJGNnpIfZPcPYW9OoId6+9jBZfr1NB6K5K8oYjhmcyTP4fGmSpvdZw+h7QlihfGpjJxrm2h
McfThgoDTuqXxxK29StZYz4MUBXS44Fgpn4JJV0Dlr9nzCvEEEUbsYfhNvPgz8URZOcvEXR288XV
PNLqXEgTEfRuS7V154iG8QifbDAMRJMQjSo5M9CnmPJWu5s3LhmkA1Q30s905irzGqbhHa+iOzKf
DDGzh28BoYTNGoOjcLyz9SQJqzTAndRJG9bbdPFCIerV26fcJg9guNwYFr7fEmxkNp3xKloO8VX9
qrIxA+vz4WuHkNHBxvRrYOkJgNDtueuN45UDxx37jITIBRk01KISelc9uipamA50aCKmMb3HgYCy
+P4GeN77+nMHbbIdjKF1vkwGzugMyvrlbKs8fadlDVgqS5sp9Q5VtWlrlBJ1sjdcsUERNBS7FIx3
HAf2cQaBjsA7Q/YlNtX777z/2QLxyw1U//KRjwvZ/Df5gta2FTtipoKjhVnmPZa56WQZiS2rYmqd
i83HY+amrlU2AhKZGFO8S7XFRdMEFfNYQBJbETmJNBnm7Zh6cmSbNyH4Tule8+7lAwH9BAb7sC6n
3gLoxYSDUjN1Ky72XQG57452lt8TlKyQNtwhtIblHq+B0HgKoDGLsywYKYSmuii83ZObEiYX5dD+
uX1hXB2UNg3cT+8bii/bdCqVi8dfqInyoOY806YQ44Oyz/MFMkqNuFiIzsk7ZVLfEph2nRzp5JQA
l3GuVZAvAF1rbhouFm5pdWmkeU2qiycdikBgqMWfN8Y2O87tN2gKGrnMj0+DbP36AH8Y3vvlY5JI
nQ/vrHqLW/c6SlWVJlMcZPVjsgR6XLQx0CBQ+H89ohSquLpC0WHcK5dW/dhm1KfPlleurxZ+MIT0
LXtk11Uc/w1frUKKPwEIT+8rZ0XPVHlkrQQN90AOMk+o8mZ8o//Ek9LXb178J+6kndN6RoDg5CUE
7TR2JYsQWQgZqXVtLGF8UV8ilgFbGoGqSmWcP5GZzXEe2OK7MPlxMoAlERBtomT4k1ev6h3ssqxK
i3jy0g38aA3lBVyhj2x/6dRuOEbqZD2rse/Z46tKxyCsYt61CYnteKAGSghpNQPfLp5Q3HOwxh0K
jk3D/1nvZ99nhvVMo4mhE1b8IutqsKXHdFv4O4q1m4fhkvgEvw7dKMweoOMid3Ur+zGSth+zGMOa
8pkD9BJab/urdrlYbkLpa0xILfBG3CUwNF96EnlCGUJ6DU4O4ZgiGi7JfN2fcVAx2ASELreOgbOS
3+DpIUNvTP0QoV/mONTI9/Ip/dhB5WzrOWdKm1qzw4fAOKIIEfrEaKHU5WDdCNQQ0dvKjw2hQULD
YeR/awNmTBGv1t8uSgWKer8CoVuDeIXICi3ZsOY9c9xajVPMYlNBov+Ib+hdhoqxrlfbi9RrVXgv
yZKbz6SNV5KFkDLcdEcykD45h9MPGcXoGWaQ+4AJHRGmRkDqkQIxGKkQYleSmCQ95JfitUJcCe17
Xm9PJ8AXvrXsfaPfthPT0+NpIgWlIhqcGahyaPNyq6O142gSYp02uJtyUj6YsMqLn/gYhwxQ7yqh
KaQh3sHZTVeXWtN70fD3XcPf/ciklsqhE4kWf2LX0EOoA70h8tom8piZkqLEUw40Z3RMCJFiWlBT
jvvA+4m0Jkj/Xcid64Vv8axYlOtSRfxRLDIt+qffrSVvBCBqJacGBTbyQUlVsRb+Is8KVjyd/lAI
e0o7Gs7bJavDEN8oPsKhnrifRQKe8AHxcJJed2Epzp7gB86uFe4QlSEpZjk6N+k/JgAGLo2ta5Da
PXGwE4ZCCPECuOXkOEpjIfEzHB+OZPFapWTB4v5IHL0AfaMMAxu4kpOUoQ/EOnLIl1dOcdH4Bhpv
g7Ni4lgLHpQp4pEPl1P9uSyI+VF8xOP5Zk4e3iUHv6WfdQuOQ7qnvPj87LVguWpjCA6D7LZdzsHQ
0kD6RR6FqoTBGM5SB0SUR39lYDPmuzv32xTvu19JXNdh5/f+y8CiQYkILqh5k6sOWPA+T6NANjPk
++zTdfoPxpAJMX4vuEi/RDKp/BHdRPvcfObUV2ofLhBu4fsFzGIJwgLcTBWl0Bmgbaqph5h96nGy
VMntjZpPhXJTi+OiAbFimA7Vhea0cRjUVubJp6FVWMoW3UC1NdVEYMhdlWiI5AeNQR1G7F/jk8qg
F+Ok/jdq/9Jp22YdiUHA84SvS+I1DBiAj+S2nYb1wpG8Ms5Dg3YiYToiVM/6rhbhxPnMWVL8BRdB
ingmsb3wRNzwAzVb3cYd5Kty5QlqJXgwahmEhN9srYTUNe+qiU0QPoAo5umS/Xi80eR2eWmVLzw1
CAxMc+FknveMdf8OQ7tZNN0vvFOHp/ZFdop9kKF5fZ7RDDvvaKnL36NMzfPskq3h2ZHRnKGv6mwO
IlNjEHla6tTJu5esAhhvCyt5tEppT+5S+CYwwiqeV/J/XRIhjJhEWg/Be+nYOeLnt98wwZUUdcNR
soOr+ZufszSIyXpbQSQ6R+uVpuL/OnmWD7MXYKzq3d9QVTT6WJkYUOI2guSYwBAPpWtsTdPe0Kht
vZ2TyX4MaXM7QtDBkJSxw6hEDvGJXY9mZ+tJGYUxO3RoNJmdf6AjMmXs38bcAWpd56vmW2+3ENxG
1b7gpOpr5QCbeCSinyLlCoAULDMCqtXPlH7q/P4hlMzRoQcJpR2ooZXUGVuYLCXfO3H9T1vI8YwJ
BJL+Rmwx79cp9N6LJMkcK2qVtlbiE0Y+MdQZrwCITIS6NQNfju+NRSBCcMQZ0HHpKEj5osmPBwYm
lglDDdljNVz4w0qpfO8IqJ01MUgkSr9vfhTn4t9OF+Qy5s2mXfWR9eoZm18ojEeF2xqUNnDAS/1u
d65+M+mMjtEZSjSlSeuppFEA9YR9QNU4Hv3mQXvAO2v42zHuy+pBAJXab5Uhfcx4LIrfiAWLBvut
VdrT1OE8arWq0fFmVPpOqNFUENDqJu0t4PmXLOy/PqanFboMgcYCdk8AMiJd1LHKfoOJUBFPvkP3
SZi2PPkeGXvk1mtTJYnXfE5iWd9CUNB8/AFBIxoKeMSLQG+nc6ZxGbSulmsTUIuF+FaoEEGKK5Lc
1yZ3LtZKZxxQgK5z8six/jK0zy5+uXwodp3Ty0rMt4h3W2oQ7ngOr9z22DIAlm43fzNIJnPIs4Aa
EFaCwwXmkPoiQpRBoXKch+HOrCHr952hp1ejBrkZ7z8sb/zUdJgkW8gB5137lrZwn5pkuV/mNeB7
/tWqDYn3oVgBYDwACEznKn6ObCQPgH8hzFAWO2yphW6UMdagzHezJ8QuUd0fWqgKTpvMvkrfXo8Y
TfwR7XTFBTZrSslPVxmQylRKhtZcMb6vDF/2asmgAdbaCWUnSd1imsNQMV/WNHDjHzeTCKffkKPu
BdA+OLOi1npUoDoxEPlEdJiHmrPx2GUnXlUNrnjIZc0rC0nA6Ae1/ShjiK9/H23/LughxtgZ8w8Y
ig9VdXA4TAFpv7ZTJQuJjI7tFE9tPzzv5aMv+9nDj5eG3AL814oVCydNmXlNIY59BWW8Ny5oC6uC
R3u69wSgcbHOu4se9NXCvWPbMJK3HkGQBqPPNqtNJg6hSoymK1lKCWsUAJyhBgSKya0sqRnuti4K
/1EJRO+mlQUjd1H+ajAT8zcoB9UZVNtzK42rB0Xt2EbePbiBJ6jD/ZlWr4yoXg4R+OZb91AI9SKX
eqa5KbaS6bEFNOCfGPXxMsBor/mJw1o75hFeFw9BD1OT5E52LvUr4JlzxdL+RbcMMA6B57G5JWBd
0jgRggxLgc6TOAab2O4uBCVjzVZ7+S79LM4iTPfIdg1nX0dPmNZWkEK6nuYUnxhQ7kqEc3sF7weH
mtlReu+g/9BDffuP+bjrjOdefwGL05aF847tlXTOyDYHVTZEP7Aj5U2R62Sl3IB2rg3OzYdE8cI9
2Uvv+pCOar+EDDGzzNVtbGe8N5SNieGMHiNNmN2MdXoohNp3tGip0crR481TET9QXU1VeNS5jNya
6SWrw9oDwTf7omLaFAc2bRZ1Wxwrqq0qj7ikaWn+680DTFZjF1pTvW1jw+1m+jWnt0hui0v8mnH8
Jz1YxrjlbYEVrlglArl3GKO4/4BVB2f7QBpMqWMkdMR30Z+CszOD/xZynSvfWSpEppzfYAap9aOs
AahXQMUm5xHiVjs9KLk1RX2SiqimlzoW4IMAQqPjvjxbKFV3qhQw9x0B4tidMS4fb/NyDrBZJuCX
yN5qgAYP13Q4lx8TZVR+0q6TkWKW3ptptA0pjNP1ypJ6bVr0E2L9Jcx/g3ecb7FuAy/v+xuMsgnj
sddwDM/YWml3UCUlPtYNhF9fs7a0/Ml3ez4Q24QHRe4E8keJItgrwb8cEBEGw2iok59E1jAtCRZX
iVO/v1MfcBE2Vv34YhaSXBciSNVSxASvT7XybHqcead7Gds5DsMRLwcGsVii+4LI7ewCsz4Ixs/W
EEcJW4XB8MNE9FCEuW1FpLkArTvVGyqOcJR3OR6kCfdeMGyqO3t9mfFSIRlnsy6BG1XtBDBd/tzN
r313jQtXFeLYILjE42UItMjQJZ5iOzzQNOi0iWQB9/C97twQAYpyf1Xzxd/jt7Ig7mHI4qDa9Iz7
kCNUa6ovPS/1TiHX7An0poq5jC/cfPmJKG1uXJJ//k3eDmBHADwTPVtxXN/jRioH7srisRslVDfV
SrCkiAKeJtCpEUHACHX2qW4bTOS7o9ar0FU7oT0ADjIiUiSzstjiUv2yCNcayyIt0tzyBTvM1zAh
s5x6WZZyquO7fn/f2z8FDSBLzrjbWelFN9oAi9Cr90Gotp23DC7LkZ8uI+Z5s0OGIjebSh3wY9Nu
5mkHD7deMexP+WQb1t26GFX31SFVfJ1XioTIRu+9NvyDgYZP7BpccUh+GRoC3bOiXp0dl92w3QmJ
/pYYGcQXRsNPbk07HPPwsYh7YsVUNRWMDLgqvBYxio0Nbme7xf7mdV0UNKGWaJGauPuij8hJQpEe
ual8pdTrkAeKxY0Pd7tJ673qcJq9X22jh+BOAPQL5p3KMa18MAotKfYxohjXkWzHA3KML2L0dNhJ
vH2TBfXWTbDnb383pPNQvJVKf3dtV39Gy/ftQPH7y8M12twW1TzHwkOBEOHqc5M+PqDFK72mqLpO
QI4BT9G+7FMW8V9dimHq5GKUHsX088C65D1Xx+9tQ2G8l6bAd24jtWGxLxaxhFmuapgWRSRxl6Cc
Y0mOzIqKZG/8XhCcK1XgTD0R8rpJAwR5AeHDcQjuEhEkF/fZx81L+GK5yU9OxqakLmqeVDcyEzut
qCclCVtOYPlx1xtBO8zyucKbpUk84FU8bw+jEPHb4XLLfzVwcUBZvF3mYoix+SK9iHkU8VBY6bs4
8U5PXBx48dgtgcdL6O1GmyKC5ewM0F9gv9w7OMvQuDQFC5q5YrmW/xbICXRmLYHqL2I7pVcOErUg
gmRVPcZ9pRBxmwghFBCIE+2xuFDN+zA6m7+XBVSHiCTZwfKbtdsz4NtuVYYOR2Y5mbvNoYmWAYRf
YAwOn8YDypW4QQdVoH2qsipfJo/NU0sPlUhIjxaIimwHSYpUmld1BMxhOUexlPRm0AuTmJFSfBNq
yddJjgyZBpLF5yoAbxv57MfGSNsKwXerlsIO6Zi3FatghmNCVgpuzUO54HmLb7MCojWrMq0JlElw
oCQGGllB1CnU/v27MnnokBMlrSxYsao0U/iCRw5ws6tg7gQreppwe3Wzuoh9KS3XdWUWgzLU57Tv
N3rkQIESoQGSoNTe6qTrirpnpm5R7u7H2wZyDdW0SSNBcfEBMPV9+IvFn1C6MJAqMJ19lBaA/r2B
5ZG3XWRVSiJyU96X3lepc/AXrm5Q/hwa+J7m8mlLakbu8/thQMQRB/IQ9ScVNfsmQh3WOJMUj/eZ
7E0vo9K/C0JstA9mD+4FP0rvDFrx/RHXyy4s4C18zSEqeUMWqzkxs34Q52U2X2xbkoWChsRWXuoD
dhLoZ0f2LrLc1/hhJxPyJggyu802xJFXmoZBHA66ERqycy7ybmp29WSUmDfprJjp8EzqDENUN0wD
BxXsUQ7oyMi10M5q104rcgSS/3j4/3Xn14Vxvniae9DMGWfQfoUB8WUXJqkMuTqfc5M3x/lCvtCj
hx5UEI8OIUHOzT84Tf78k8v5zNdo8zRaoziWDBmhgUsxVxpUX0mPQSWULaQVRDwg4Yq9Lf/ga3KY
NPKqBZ/5pZr7ICVrW6aozkEfAX8UzLdIqoMZbsndKVCpEl09+E1MWgAMGn6GZa7xk0gDJ0uy5p9Y
kZjLdhdG0uz9fM2KIP3N0/+b2qXbHuQ4QGkNB6cwOcc/Hn5T3Tu4zpkgRc/IfPii5Xl3R96I1ch0
XI/ij+TGhmVk+kldiwWojopqDtbvRGzLxpVbHBrTUHGyxnl3c5AJUbi4Uwu5eLWX16/1aFbNkxWh
VRGICT9A0yT8L6fIB5nUy+a9dcCFnqOG1ihgAAceZwI5yEa0yZneaX02IgaWESInpzBXwq8y8JM3
GzDt/sShcJE88D6GQBBop0oA7sxHHo3YjJ2kW7sodH9//+ccdknVmJU+j1m60NYbgAsqCU6BPPWf
Xcl7o3pXLAgC+gLzOGXlmIICPXfLocgqPKeFsEq+tfxFCqGoGJ5FI424ova7T0OQtEWmoXH0IWAZ
gsbr/QTDnio4sk6XNJJ7pM1Xh0AgmOl52G12GiK41Esv70sFozNwYe1/+wLuqJLmWD3mEwHT+VXC
r0o6h9o0kwEsNJib8BZzUUDPwfjpz5Y/2x30tZ+z1hjIk4sod068+KaqyiWiSDfAiCNKjoC22oy1
3C1T9m5li5Be9QWopf8AmgjCH3TtumUlTd6lR9t9UHvX42LoRceG3Tvm1/C6Hna5l2nzw+7IKZNS
+Eue89J94D36kom20aDBwEHDO6k5vCAlo1UNr66IjhJ4WkELosiHYX6y8auHsEYQsB0cdgWgU3/z
cp93lY3NgM2a3beo3QdrB9JR5gMsmXzDd0UaLBB1nk3qkf14pVB2yHfdVPnnYl01HkLqcvb0kCXb
E0wBADbzH9ZKHaINMftB08KaB7m2HZgSxT5jCGV1cqCK6DmaHy8tX/7vMyAdIBn5nBUZKsmVM7sD
zyMbANYl0i2FcWLtWLxHg49ZoOw/qRwpAtxcj3ecELcmVXJDqrRLTZ1nNcCQfudtgfWtvo3IxCjT
PH8sJQGMlAyiMEuaO76+XlmmTPEPpwcgmOHKTeumF1FsfBzRCrtpX0JbR9pkH3gf7THMsCjfjvs5
hAP4PVyEwrXhR9mtc/+u4TUQk7qWDZibkeWGq79VjCwQq4vRy6gWBdDUkEd8GttOuYOIJIKIq+0t
wofEwYG8wPfOm4/5RrGWGoxO9/gYDNZQ0eFfHTlDMlcjtekx1zqrUhtQ7VA1zoL9T6j9wy2Gn6vh
krvd/b2vxDAKCz4/CEBh/MYiHEeu4dfYjR+ZVIxXlOmG35Ar3eEJaCnu2LRLi83y6Y2jNL5hETVF
3XKs2jaUPioFPHErlfSJGOsiKZkDRis/U+z55Z7fOG9ToyGO9k5eXnQePqkjF3tVs7ta3AWcaJwJ
ngESW6EWy2WM94QrnyhgUyCtt3CPd9HmOr0SKbE4z0ov5r1Wv6Dd6tjSqq4p5udY5bOaZA0n6Z07
xAId3iCtWUFxwpzoUGmjE2xWT+K/1ShQXxBtDRQJgPIoHraxoYWEgVi0GmMXQHltjkl+p+fY9H0p
mUWudGsJJrY6/KqDjqdfj5hVA4PGnZzyw4GsAi2kInEfCPSWTRgulczQZu9geOQzr/4XJit3+Z/k
U+f6PZ8eexbb8cPYrIW+ZKvSH/C6Ig3K41qFLQqTtFUgAePCAzGap/iHSC5YYkstPiYw+4QY/vLe
4i79GjtpN2GZ1ebaOygtvIVbDSvb/wdznb76dqo6ITE1WLq7MHfnTy3NFDprLx9vTPmUdzyPBuKD
IYU93axr2xJa0Eb2KzVJfv/a0GIFf3fef6+bFQKj6aZZlG3LKB+9qL/iduBQAXe+gIs2dyl8Ylt5
bhl+vU2WaJNvT5se2glo8YOoI98avxjthtqGrJlbsWIAjtO2k6iOwte/PMPfat5KbfCL7ZE+NqdM
Fc1e57YSs8iQv66XuXrY8ITYmFYwdBQzQ19QwnfnXCYMBxpLGB4Vnljld55h6GcMa/BJ8CwgIOMM
RlGDQGyNya8zf9zlR3kMhvzrgXw3iHbatgQQu7aUQ+9CksFCq1ha4BLpi4Cwn0N9JzdoKF+SRytd
AmEKa35ZdrIOrslKS+31h3GotnsMs9gUnkWSuZ/eBwXmv4fElhL4tyLEEvxUZ/Nlq/NpRziKuiz0
rlSSx4Ui0AZt2aV+gDUrlGDwAx3A8xXaNdju2X0xQlN558nntR4Elt2+du8pfNI3624A3jZaZsiS
g0StV2VL/YUemia8YuZZG5LSfBqU0SkdNo/A+j7xOIrqWOUA2gi8E/vbS84oCVdbZdMf5++gqOUn
gWKEgTBy3R+ImX13LmCHrAkYjSS+eUF/63HeMvgevov22Vu/SrIYQjtRN1FrnUozVWq2KduyQovc
shpkBg7k5ovQYO7E2u4dis37hCq6xK3VtUxKUPoYdLb6uMH1DzpMJ7H3cZPIndPgLHcu5G7hY6IK
m8wUwrHMmE9FiuY8QXFOYiyYhA7dWVrVKZRryx//l+jjPUJq4pLsur7WBn8lDmPr11Wv8Gm77Ibc
gGGK6XjCNB4cT0Fp4M6mLTX6u2/hOQZLwUb9QWdV5STLhw3dhJw4L6kosZh6m6xxsScJe0bgwGqV
ONZrMISW32nYlUi1yEgC0447cKKfv2IL1idzkRkDVpveZnyb/IzGMH6MeLRlbf/5I9j/8GqYYKIC
UvhRXm/pT2DHjLW+zN3pNgviR97C2lMfLFK3iINjbkSO7c41DKo4mVm+Lpn40a/2SyWk2ZChdXoH
a8W2tVSJxiEtjJGixfI0COS9qRuHXS6dO0jghvPFEUfHA9ui+1V7zwyFCsr6Sd4ntvdWvWx/1ge0
S5iQWrQiR0IratfpjWtdBXGmDS4A850lqLBbH941+0vm8fl/B1fMtWRjFSy5UJB2C8iKLR5+yfEe
7HOyQfM10P4l80EW9bNtZjxaWQxYL2AHSAkOdNWbvg8eg7P7cXU1PC2F5nmYJmR3QIDZm/dszwuW
36hzLytQ8iv1ePb7zMSpLUT59h7rz7xN/CBrCRq8DWSXH7ly/tgOqZoXl6gnfcs1eXhRP2LQBDdJ
kN1bN8Fnp/WHHuG3r6fp57r8P3vAmY5LJOWoZHt7ZhFCzRE0rX7kHM8piPTL2hRQb2pVbYT6Wo6S
zZDsuFUiOdz5l9cR53Si1sL3Ynp6pklX6xY6/X8FxZqujTTFkuXYuGUS3KwHACA8qv+M3yJ6eVUu
T2jvcn4zjnNCh13wM5IFH3eL1BbPVONU9s3s69tUkoxYca5+n0EzyvYLj29o/tx3Jn5U8c5pzq98
cBz9vHRWFcuCtmOHrLuqzcfKkkS1w+8NpPo0OZaIHQmnlwcwR63OvlASvnYzcCgu3AcJ3zc7kyzT
G99HJItb1qvrQcg96vVjIH5CkDr7y3/lozSMaFhwldI0S1nUujMeGKzWw5B3ubUPcdPCH0+uQ8hl
vufLkxciXhVJ1/rOIjeU8yFoMCUMQTBM+AxVW4KPOgg3KJg5IDB6rmvY+MCGYnqjyUSKgBNWYZpQ
UreWoNmzW246DxwTXiockHpDvVBPMXi+rm4R5vX5tYOjMU6CF3uWkzHNNfDxIJ+LPiaAudgGQGYT
eALouAaefHshDHLjOrVmda78dqh9a4vVBwlrpK089lieiJdZlUil1fzosfXB6UDD32DEhPGf6t+x
L5wt56ihpnOAKkw7+dbqNqBGizQj2yk8elbrXs0sBrR+QRT5yYNOzWMHMza7sMh4/FdKjQ2ybO1d
svqfkn+3NVHkG5It0/UxDKmMOOABf1/sfwgzXtJHiqa3NsFjrZWV9R3B18PtuheqIrxzWkDQc6Rs
98Vt7X1eBubRsg04PQmgAMkVJtPROYZzfDj9JQO0mhMdP4taYXvCVZOZjJxjmoxeh5ppNiFCQgTm
k5zB+DUwUjJxhKADM9ecNH3YGUgSNZxQVJT5+POJ8R2XATOX7nxe/j4sU2FqtGnt+GwbN4rdlw8Z
K9WE3FuKIvd0PwuOi3/szaWdl6Dce0/nqkTVQCrRx6S8YUoHroaHQtKnLwGpjcz4MqqfUTweAHsL
qf+4l/m+Yva75Gbdn8PX7ea6G8p91rRKW8SPvQt6jyQjRd5bNRbWmpBnY4gTPNrJJCqI+5DbmzTd
HI18BRe/MDKlMaSW5mRUA6JFBp3nbIMOshsWWPWpreA+Uhdf5cOcwBjpwRVi6BSw1tuf79tbuKt/
15FktL0iSRRknX3mqV6mQJtGypv3szo3bwbO77t6hxTOwBUIzVfH+UvWVSVuMonR/ACI4wpL0gHQ
6VmIp8eDKXhhBb8XJblGPEheWLixRpn1poS2PXxKTYzj/s34UMy5A6ynHB7XS10tc5G3/fbDhjSD
yyHUmMrWtqkpZL4Jpp59DVi07XyzNLqn7T4dGHUIv7yCtzwxlM7hePLj+DsANK9aZomNRdvZ3l1v
0nGvHfds1JeXbpx98DB67I3aNMuSzl0Mchgy7PrHRrsNZYy2I1WW4hG0Q0aBZLoEjcoLjBYdjiY+
6PkL1KQjMsHqyZDGW8fsOQBBULlmLlV+6KD3aFugHCWC5zIkU7/HUf/5ER9D+/T3ixWklNoKKy30
r/9LlQr6Rz09fsQzM9CQskND8aYPoKnm5x7YD53JKY1VAdlBXUhz/vKzMuQYC/LbibLF0QCMoLJc
wheynwXWYpeK7zpAAZjdqk18h32CPSOs+D+9XBPaxjJlzaYoKTCLViccsKOTVIhvH8OAxO5pxGqO
IvXuCSZRnON2HMABkjfHd9mVRXQnnBh6rDq0uYHL63J9af4BMaq911PkOLj8USW3o/0DCke8kmTQ
eznKjy1fTukwydvUT6jT1eo/KE/nvmjPjxRGm1+Zs3CF1DPe5jP0OnEf8nlxCikmrH9XdroMgK/4
rT/DXrZevmUSvIr4KIkRV+IbDXdmSywvPcure3PNdyaCFwYAyiEyYyf1qd0T4RcmO5eBrxvspAHI
G7OtLrCkE1SCenA+G+nX8ejL4RHUNL3IRcNJd3QOuDcqJ2g7V1Z9X126JEYFRa2lwad+HofhdUgU
7OOUCgkZxlVU+c/N1qgeXr0yPyXdoPj0SY/EcZghF7I0zj3/ZG8NZJh74rMz6kooqWWacCEZuRvr
e706dxsQaLiDJe3Xk2G25T0/K/X+fNgQn+2ygcTkwywM4PtGjj2wGRQU4g10U/zjrOQhZ2ur707I
7utxRRe9qXt2ZMLRuHiqXjF5lek5rXVGzVrHAqLu7k2ZoEtleY7TReI6YGHRY6vxm7wLSMZOpy6c
kbolC1BUUAB9mbW3a30iHfK4YtkI1Ld/owyNtlc4Yn22/rpHbl3JZsm/6yAW2n2+uZnnBGhfWB1x
kCAy4Uamg+I+rH0Ml3FS7QlMj+Wdbz4qJ5+DNdQTeQLNS3q6lYT7V7eZAFhC80/DsD/YKvop4nQV
8wiov2P3NmcZ2pe1AGNrYehTzkIBA+MI888yBMhdEOlOGM//xgjqg9JtS9r1cgnJts93WHkI7Tjl
qBjR/oABxCulF6YVjsuvpePau/e29OcqHMQol1uS/42GxITncBqVBXQ3qTT1i5oug3O3VgpXm57B
eKqbm5WJu1xhIeX7gddbB+prvWSOgNMqR0aKxYizbTkECrYaxV3pD3XZOv+R7Zlm4c5lVSunN614
n0mNhWCAZupyD4jXqTNFNeZKTARFBsmCGTwRB6WTNKYmM2aA1fPHicNdAxQjMaYqnoVChwt8om/e
ETv1gfuYYVuEFHLzik1SVHZMcOlbeJwKKobXsKED+/cFHMPUvlAlwrpicwpBTAjjK5SGtC/FY4Pv
vhw+kdlquwBD8GKrVHAf17T01UpCClYYKkF1u0YVSHa9m+YspfaUxAcD4gTtullA3s7ySOBHNN5m
iaYClxkNjLrcNMsFDxiC6m+dtoLAz3m+XlzeH2GCFJKF+3CHc6sZbSDwrfwp5nlFUDpav/TVg02W
Kv1TXEtCQfgVwa6D66c9tgN5uw4yKCU3TGRbXb/MnJyILu/WYgQhGrCkzwxlInV7Ev2TE3UWeUaV
fuSOuKlG0NTmD8nYQ7RFqpyLyB6DT0lDdY3luVHayJKUGSVdHsaHJtFPhY5aSuJPTCQRvaOCKQVh
o6U1GD9WWtKDyXGGiMIt47Z8m25iafWC283aRwU1j3HgWDIbmDqM5ixfRj9EvcdjmNtUFm1QreZq
WwOBZ97sUgyVHyNhtnBKkfCKtLeWDcPrwvXK0DRrrdh0qiVc6o16/yvQwbE0zbo2siAlDIw90HVG
tbJUuog8PEdDXdN1skjU8WclWN4DM0x5iZ4v8iVfCxhzIxLlc9EdqZ0ACV14reefEvo40JpKoNVE
MNWy3wsT9OjsFUs1NAs33Hkgl/Ofq6TaOQaGGnUuknxgRUFzo7O+5HxXmvUPi+kZUTUbzTHK7DJ4
1L0vrGGhpmqlzOPdiWmTiMRyFhBdxVq5dCtAoDrhvPL64da52dNskoMRWZMml/OaYca6jeEZ37Ea
p8t4djHfe+RDKjtruqFofq3uI6V9g+on/1umYunhy0hQvcCYx1gixsMOO/342BEnsZ7777MR6x2g
CSSuw20/bhluQaydSYiAM6S92pWHbMUhWiIu+vkNGzd6DsAc01FVkvDnKeqmFNIvWrk9umuGN5qz
4yzIv/73XxLzZCDX7DmHCGJDYDAo+AdVUXDr4mL5ACnhfnuDhp/l2AsObMhZvynbBZo4doBrGwbm
ISuzJSci2wkm28Q0gIHSLfkiIPT3ofzh+Fz8SwGYh0w9grAYADbKuo7r9qJo+tI8NPcyqfBFym9+
axZN961JX4zetapwDLHOaScySttkgUN12ujAouoyHp4yGCuX6djWvtuLgPOD5LVSv3hb2LGWpkjY
9AgG3getyg1A3xSeI4FGX74/KQ812zx/f6XuSy7Hd+K3ulOas3K7UrPbjskxcKQhpz7i9NoFCtfG
exxUq55eIpbuEYNvB/GIzIlitve6udqaH4zCBec5KhG82tIKXaOLAJwq2Evk/r9FeQGKJYW7l3iX
/1Blfw5UJ1c6zG9uPTyoPaiPNBGHBDhXZbhvUR10foyoy5sXTvyzcp/wRZ169Z05Bb7qiMZ/4gDO
K9A8Y+iBr5wFmcwSB5KpvcD89gNSsZ/xsKcirLe05BiRVqdWICXWDG8hRxuBNK9DTNgWYAw+J0oe
i/Sxxg/MjFeyu19vNCB6pv26RRJgk63rsz5RNTLzhU15/YPu21Yg/f1Jz2m0d8N3KdxAoDgDaPbN
v+STUXmHr1GQ8hL9RvSMSS+H5XF7lvMgJ8hBpE740KGRkvLnDinuh6yWN0EMJwPrjmznirxnTCyJ
EYRufrRVnu+QXOOMmw+DRTdXqWGgf5pEprWpKP4M519PbJyqm4Q1Y+gtFMB6QgSVw07U5opRefF9
mYSer8urTtVWUebbHlFPMxG5DH1SvJy4ey0CM1lkw1MBuNPugE1UCySR33vEjrBoBLIE3RU/mQP7
ZTprxXEEc6KzGSQdxmR+YzBIQD80tIMs4xeoh/fVIN08pMfP2s0XD6QR6Zfb9TvyBDgNJmLCyeyB
DGH6nxqB5m7qlx/KL7ks65xXQjm7in4u0ud8bz/VpPF/+deDTIf0ltyW6HorX2hW/IDuSEy91Rt0
avqyQDsQAWCida6VU+7Znsi+LWx4sYwEwXEzcg9TScgbbxL7X0mKMOJBQ5DsCMiL6g3GqBwGmpQj
tp9fqWrwTN/AXCgwr328aypql7Fe8Oxp+ghnbMbLSpYvfYtJKiLY9NwyGczxgkYx2rjV+3xLWrkE
tWlPrL2PU7MiliI3skNegn03NPhFgzsKApuh4Vf3skjKkEAbgZX+Qzykr+3Oan2lYqgeMVpFNtQz
0SNADP4g6MazHfnIVrDzfT0IefP7tWSK/0QnGLmNJvCyBszzD+bwDMBMasTEtJbZtGz8RaM4r7Yx
hi+WoYA+Ms1SnIPWO8Fnz+WKA5DhCi918lMldZsl/IjPxeOeyL8Ac64OW2nx0jkcJ1cbRKiXKNBH
qq2RkNwNycVpp4VumqSNpnTKL9QYq1aCqgXceCT/t05ZmfqR3Ux4Q8uPM2ej5JVzkKodA0F5Ov7C
sf5hEGwHedv77wjVQU+oXf01ppoUjWI9eLtn5nSaRo8h96KzDXGUJD2gffFmtd1jIhj6A/1NvP57
u8MdeS/KFcRZm1GBN0jrRxNr598KEWNaq0cVHbMxcEaNVC33pYhrodMN0IlkqDJdBXRYzZK7GcrN
eo/d4Ur2hM2uBY8j2j93QsbfW6u+64a8KtybOA4RNhPlFl7uRdAiMI4YDmiWov6v1HKkZfLEkzfH
Wtq+WLffClri/wcVHWX1bHDdfksn9YKC9lTYMSSQxjFUQgBTfFLIIaQbfFggqWoWxaVkh5GLExBL
+pnbUvbU40XEIh8g/HRdseGeY07XmD2RerwnFbf/QQA28GNnVk+I9DSWWALtlnpLE4CwH//krv4V
gMdmjkkJmmv5voj9UVvfRuq1CT6N81NAsTakIDFrB2j7MeCWGdBi0JcbN1Ygal9+ccCYhkDsa1N+
lf+5bHVIsn55U7WppQBvjiGFgTnBR6cz+PaMhNroujsPaoghuS7fsTpUSHogELGEbD4OmV5ckTMo
cwjJL1uDJZXpKi9JW3WaqUvizUgNaxCQdodXjOkJMbiLfiTlFKW4qOvSjooa4r3RtAhlQFXL7scx
zv85SsC3zGI0sVMwaFBi3L13jMzVMJ1OPXy+Zebo73UJCuGoUQWfjkURrWsZERW2IDGA7Oghc4ny
dDQKKqfEGAEb6F3ORHQgUsdWpO2DfzzganIhJ+B7dJ83CLhrd3jorXy76exrHdqr/4JBzoPJzr8G
oIr9Tw5Q/VgtVVA9gBP7QbE1s1zGrGSCCjgq2CtA3/2e8VxEqeIs7dfZvD9vk/5JaF9AmYtNAoGu
xm8F3mNw+p1h2J7GvroH+TteY33U2ZGJf2IGQbsHSDU+lrrBjHzWOcBsaKz+QQZqBRZKcr9phxXM
X5v6/cFUWqbhRkFIh5KTRXMWCIyvErdxqBUKHe7z+kj2/pYzh9THh/L+7xSxgdJcZRJQ03c1f+cG
0mW5MAKGHiW+F+j/pYahhN52G4+CBa0Hx8pmKe7kAqPx7YwRkXlQatpmqUEfNDL1vYkEN5hRbq17
BxyocS7Ag0vAf5E9uqBxLjrQQSAaIcDZWtzSlqBoa8nFgsiVqO9MV0/4uda/mYlmhZdsw6zkMjcg
JCaFGXRUlTAn+tNK7digNYvgtT+F+Sulsvz9e4Mr9mv7Ynud/M+fQ1eUYYlnaqQksXwSflXou30C
A5qsFCRUCbPhS24pZXectPLC/pjN00jVERZs1LY9TqWOfLn2Vi3GpzQh/vbFOJTbtL67qeVSj0Gy
RkG0e6lvvUUqshW+gR5JwB+DLpyXXLTuc6L0c/z5m/fXpGg6mXI6qCTHB+pULxrvh2qnFh7F7jr/
jsNPzNKkRFmIQzyUOPHMuYp4LXGz9h7kgh+auK/ML4twGPxEdxnKCqBqJMzxHhbc+GX0o+3g78pj
6Nsj+RGqYwWmpWFDWuSwhA1UPthUsuujNlDrZ17fL78zwLpyDmlaFNKwHgOK6sHPFxOkoPgOSYlD
6/P/u0FK5ojzSejUX7zXn27NSbWP69lrPiUPJg2Rs/R4YGghPndnJPn4HYb5Q3gGEHY2WTA6EcMv
q8klqXvv4A9fAKnOCIduwDEu3IW47r76vyUeIFUo3JrkUWSQ6RUcFDKeuUfpwqFIZI8YcZJP2r3k
NQjJB6Dqwj6y+daphQLwNMFGcjEGT5ZhBDrO0OgVEQBJY71058Wphbt9SpXTqORUVNk6bMDtA9gS
kTtHgeJ5bOPmsfzYtY/S8SbuhaT0VMmuz/WnvhL4kNX/qdphqfA2jM/J2QbqEFvvpnu30LnX0ppm
TpvvwcBQGbWPTHa/DtrxOYBZ853F/8ab2+5qSqREVS18twvqDYlWhGvv7/Dcx0NAXJpkyPntDnfT
dNg92Ex2QCWZ23Tb/U9wATZHnpP88XjTo3nNERnf3eMZAvOxj9LP3nlEOuuLDYUWsY1RhY+8vgHq
Mqvp9fmcxPj0NOUxQJK3b90aFLznD66mHYfI/05OwlDn4uojGoODBaUl//+B14AHtAhvPzYhPbwc
ooPTJYEm1t0Dqjctf9lc924QtY/PhhKLIQXltpBwxEPDC75szlEWWT6tTkLXhryzAjuqq3TJYe3o
ITLi5bzmIzsUs7Bta46QTm0uuCIxrFPZA4Z5QfS3oA2m5PY8BSWjp6XHTfhiK1UtrbP3r0YvOyxJ
OLUVtDZBZhNjKa9rYjfGbJRydFG9/3So7N2PZEjqzbIcl5iqMF5k3BQhHxZsPmvHe89CDUZzwDDX
I3DoEkGJk/u9Pjk9Pxu1DLyf23ktrWmSYLWfa64X9PwSqrnSTyYk+EKKRYplXkZIKWN5ERy+vo9i
BG+VS3fAdyE7jZXuItKObaHTWVt5iOy8Rf8VETcQJnbwu7XhaYoKEeuwufzy3OGxLLKegvwBxTpE
wRyUg4vlGoBSpM3vT0GPRE2WcdE63lBpRug7UtT7iTaz8oeyi+goaHjaaIK5de78c9I+X18mHDqz
BW3dSM2CnVCYngwXolISqhFZvr/2Q85VDOLGbQuRAWPgmKnyy58zDAN6omTCMiQCBOiJbd1ZozRu
kSR7cYhItvo67QTl6S8c4f+v1FFrpQgOEXLEjYktAgujzgrv/Mtdf4tBoeQ6S6oaDqr1bCWnkxJ/
cgcM8UjywM3J8pbafgAmxqKqN5Je5g61mqEZm67qF1zbauhsQ+7KRMSx+rNCuLwQ9jZ+dDeEHWbn
SX5/cPi+AujWpBk07Vt9Zirb5KHqiXKavOWty5SlS3naQaQx6/IJYvo5DJ2zRozQTjKY7MjFtkd+
wdqQZHzTG6WzQ7ang9jNheu40qcmqt+lFMFO97dJZIVmlG8BQvyE41NlRditpBGLpLLH9WUPrXW5
5VmYCFhb6m85asfKrHuxpnD3gGdqvTWSJw5wlQsORPxzGpsoxfoV786Y6PNbGrjkQJDAAoQlpAA3
cBdVT6synniVO0XWqJ/VeBaUEQgG7RAc/HsblfIPoePWnHPTzAqXFaHG0GXFWd7yn2LZscY8ahLM
AHT7BNfYQS9lLJA8MCbITcx3w/lZ1htqlBbSgwafm2SpHnM/eDBWLGOX6obGlGGcmezRjXsq69kL
8SJF1oo/3cMUdRGelMUP0pQh1RKNjhC+ZUoN8GhiAlPVIM0higMPUZz+VwpO8ctW6juuOyqRk1qm
9WTkIyJ9SxBV0d/L9iMVUvXCwZHFehdiEkviirzEcvLMc0NmpGKfcw5Xd9sQBabBfpTKrAV0IrfR
CQcKGxnexdC9GhJj6ckCGND8X39s0h68KONxeuqVUUwmiQppeQE08//kFm7KRgvqu8y9dw6hNh/Z
FeSydxjvxZms3GXNMx7eDxaATEvbGQqBQxt6vrgw95mApjKFXhD2v0MZj88i5JkwknVu6towO5C5
OiM5C1+y03s2ulCy5j+pKWurO94Ir5K+VMeBT3C0WeBRaYPEOqwO+zhQsZ4uGEZAOIoosLdvGeRx
SwdJ43INb8DOu9TY83VursQyrZBjY6UBDJbdPY6tFLwVl51q/t3XpL3fKzLhiA7oe+ra7C1kgW7u
BOsY501gIY1v1QJxqHe+Dm0SYRVJs8VHRg/mtkhKjC7kVMd0I+/BkBvWbmGAtAbJF0y5IA2pkMlv
I67mSpxZg50aDtPZ3CS6sAsTbWoNPhDm3viIV8N1hO8RqlbAG73qRqW83Ru8XHF0mcUZ+yx+sNqa
WoenWZK55TMAWJtODoaHs9enDJ9OiO0W4KZYv8Z5bnkrvzwaZi2gd00iM85xHz1VeYeUIsXdMJhT
HRBAIbHVCXYBN3tJTmJyf0YZgjFybQ8hXvYqx2czzVWMLlecfoKrZ28k3kC3Rg3HGnJCjO8BxLH8
Mj8U5yK9owePFI4eEvApAVI3yQ1h5+5uBbDF+j1c9imuVcCL/043aPU37HLzhk+3b2+t1mZK4mP8
udN6W9/1OK8PPmRzbrmNGwpK0OnlZmVb7uEKj9gqqqdI6DAc0xjbzBXsqk6pEOtNUKQ5yTgsZGON
seTcTsZIYM4rG6DCvqvS8m1UIeBHmh2FXeqGORtsj8rVRBemsJJE7eVaxPKsudmPw+k56JiA7ic3
MhlFMprBQy+lSOfd9J159E/BYff/pxWI04kUfZt8HUzNZA+RL9r6DFdjlWKhW4XzR9twp7wB91L5
K8AiT5SrtbRe3RUs9N0ncDogbixN2EFp7Jeg9F3JF9ZDEAsRAjhMDy3LvgO0pv/1uj18Ed6IJqMe
lc03Ceg2OiwqAkft85BZYx4TOzDuklh0NNSuWjXh7R0PgW9HyrA+pU1w3X3+gjZW6AjyAOMi6lbR
TVsoeTavzGe5Y9iwLGJRcB9Vq4XS+q5pJVBvk1mAik6mGNzJvSUSPf5edYJrkC0fT3JgwxL2UMbb
upnzZGZp5owenIfFoUjj8WZ+tnXd/W772DLUjIZ4EU8R7tuV83DvE/y+ZJs+2JdN2N84wclX8uu2
F8JSW9QuQoHXRBbmKwzn2dvG8jU+WCnz6vOFVN9wpR38Zgyate6gTfMpLcxag2FJ3zAjbrGVnKyc
0W++Y2gKXLOpTQDah3vOoZOVm9OEKd4vmcno1wQiM2d2oWB/+qyZoSBidme+tnL1D3FquQ78AVgL
KePpXc2bWQuHRrafMn4xifdhi6r7aFfSiT9SgSGQEjb5eLD3FCZYzb0zH0O8WfrfeK74r0eN1HsE
VYZ2VbMwWI4iSnPnFFTowNBIUPPZF9E+LGn2rQeVapsmjcshx9uxBnoJFkS8FN8kGVLrsdvocAkh
3COdmSgVOR00xnm4WVtQCMCjGNbkE9LAiDsXSsAbSfSnzC8la4gpzc3QeTZwUIw0VLDQdMayxFtU
jBPu8zk/rAy1MkP3LuRzK/9V2qbMLnULurPqM0t+vGCmZg7KTMmHhL1fh8l1kdBObxARKJU7/StT
r/GhMxU3rE/3Rusyjn0oMC9YldgWmefGFW+nfgzgh7kKUGCkbXJYpcWD07IqYL+JSULsZFn4SYCc
hwsPhDDng3FFrpXjQMsLXpm66H+hFucZECpXJHiFKClBwCW8SrWsFuMwDMvs/LIscowBT8M0DA9z
+J9WsOKNHYWBtBqUiklzzuuXU6gEF1aqkISg9mHHs7uKCBFlCu92Vai12vRbeLrEfsL64yyHzoLr
6rAUN++ZQTIWPKNq9qgThs8SyVo40TE3j0IVhnOJrhNBtJj2sw9ddFd2SE3490I1u9VQ9/M1CKfg
Rp1rxCS4wtAy0WpnE7nAIAO+Pp+gn1x6Uytaf2Lh1IwNxQgqp5kqnNiACIZwM370c53SsK8htqAP
KZVgzE6cmEHjbV3F24jHRI5yvOmiauAYApMoO/KXD+vkxQcVOGJJX2Xwsh+YQYx+Nb+h3LwJJ+ou
rnb0JKdqS60vOcGUoyDyp20dvsHqqLjc/u9nCSUbyzySCU0DZI0VSXdRlXc/06cM9p0bEE81hWyA
0lmdDCerW2cNzx1mYDWsMxxsEndNdNNGGttUPOWV5KXEXq17XqGmS8CnG7A0rffPRvXFjtPcxnCW
5d0DrEyIsH6GVLmGBRGpmE/YTZ9S1VVqpJXkHblLFsBc9o9+69E/lvNK4yyFPhuimqg7f09YDFwv
sz0SpIpBYgw6+K3DhA1Wpw4ovNhJuA8ZFWBN8SogUUIGXqxLcNJW3CrAgBlkwSuU/i7NnN1dn9TX
DngQSn4iTPR7liK2qRAKBesiW+CGmY7MOO76VhdmLAZglDpJmOTvuY7EP7jI9Q/hFbt9r1sZPDs8
kmuKH8etoh5pHmvV2YXSDZu0YYtyDOmJcLmUGDND7y6WBUjnqp7fYov47d0syqi2Pz0gp2aGmLg+
Co/ds84TYC7uWiLztwPAYlCHkU4RIy9GRIoulPCrD3M8JTchzcUsapFIound96OYun7ezkKVY/qt
r0TQIWBmj8tPc37G60Jj+DVukr5Q9gA69b5oowtE+wV6ESiTEDsD9dP7M15nKFgc2cNsrsxSw6zg
ntatLm/ktxwAcNPZDrVdmeC+qBGV0ig7mo6GBbWJq4ZRqqn+596x/a54fiMzMcNb1DkI+Pb6q8x+
zqrbLKwVdSBiZu3x8eqhMQcZYQWwbeUFTkRvPT3L3xtDOH34yaNVzaPTr6XUrNsNimrVi9KYBmp5
8xWlUDuA+gjMEs/WSjRofNHOKuWMn0c9suFVQxS6iLHwOtr1DWtGMCYZ/ekHowDpLLZxVi20i72l
PZPjrM94J6+ZsMp5dRzGwReClu8+aqrVdfCd6ta7osEC0k6GLGRYjEtUa1u7PMHsNtcz5S6fn+KL
LrzSRCgDVvGgjVP8uXffCbAUhtNxorocXeLbL2yK0cPrlrldRwMsO8W7BNByjm8/CU5pNmHv/2Gh
2PSnZ8TCaiASaRJd8fNcvNgjtuFhD4vM9JgtaYg9j1UzGheDdKx7Rg3HjdMXtf4IoScMZoXGpm81
UgqW3DdIIZyg8f3db08V9YQhPTAguXM1mTK0TVDL4U+qnYqUXe3Z6KGFwGIpLBgYwqu2Xnth28PD
Da+NQgUeRGG+JAsr1kB5eoOmxTepaVd8GX61kR1c7mPQ7wK1r3tQn60iryHX7q7NvEkYPGlkYBzV
v9fAGxAeWoSLTXarIjCIS7yb5yymFbzlfniWSvh8W4yD244Wv55gUE3ZQwoC7tONr1HpYw1j8uay
UiPI8OuReck6FpBOxHsFVGxsTFJZnkRRjHlHIWRKoIS34y34Ib0INBnwNW6uP+89WeO+geg32m5X
RxhuEdnArqalP6TizpfZzfqT1W8C17xqmpSxea6ONBB+h/PVTVMQdzRym7cY279c6vjhEwN/Y+99
tkiQ2w5o1H+SkivuPZ5NZOOtuxAiPR5q0M/veJxqpQ7PSjgTJXJ3gPKQUwAki7u9B7juiyA5Pv7+
/5Xq6dL8LZShc0Zj2f2qO3QarThb4ywltr7jdSgfTCE65WXQ26xiX+5o0zeeaHWV93mW7mbILXgL
sB3X92YlB4TpLleNyKUioC2JvvNYu/cEjULmMgR7xb3aK5PKl/Qp7oxdCvbbzkVfiJXDoaZ2ZfVm
mEWBB02ISxXcmmLEEkh5M0eatBk5YG0b2+IPLiYBJLf4FZluGFAZ0sYjDTuHxg+QxAHWwz6FT9N4
4P9HU1JHz3KWsutZeEyujl/zBPjB23Aq+UeVyYNZMmniTB74l8WUE7OTmUWE0lG0Lbvm6pj4KMVf
E459Jc0Lxuu0bRXvQPbKNsmsZ+EAEBH6fNaguHIcICg+f70MBUp53ALrb3SK9ihRNZO24ZobwX3H
ClhmzHMb8KwCSW5e+slDpTgNVr01kYDgCGLwcNR42/dGJ2DjGVTg5vu+TulxCmxTFBUM8ofgTalA
qk7i40mP5Z9USepi9I8aIB5LvEjr/16CTUaMzgWkbf7Vdunn0nbueW+wvCFz3D53gWzPtpiGxla4
m5p0I8LTtHBAdmm3302gjVSUPFPfJd5s2Z9PZW7qhUkZKw9/Iwd2KfwBJlGtk6PmnhfPFYCizgNX
N+6CFeWe+Ctq/MuycCAYGT3zey+hok3bfU2JwOva4LnC+obfCkfqIuTynj5MQGPSlwipUx2o5VVS
xhJY+/4xDXYPpGK5qBz1f9PkR4dIYp+j8c6gA8Nqe8sds/ikMRofFUbV72gdEimaBW5Phk8PYzVI
onhkmJ3E/HcNv76L/51uwBJdZjx4B/hGpyTzeTBkFDQaCqCdSzvFDN8arI42yEX5N2N/NdkNu/yS
UQ+fpfELk9yNpLn9DB4+F+w85WwZmWShO61U4ohXDGGKHRw4tES/oxP7OQ8zpxxPBIgMfwJu0Fx9
Wii3aeLjlmTVG59C8xpMETDnWWwvVyvbnU/QudWVYh04hnK1RDmZcnwslgM0vJLTmeVFv1A6mhtt
RM8i3ifF9FcIcmSyxTXWuxhoL7u32RGjPyQwlG9wVkEyiwHKJObQOqj6yafeOYEZLFstK0ShBxm3
QxnRDEDyp5cQ1clCjX1JcHakpPKZjkwBGBzJKuD2PMG7tSQIX3LupVgLLBK00IOCsSp76/ietsN9
PqSryHQ5kowtbAAW1Iz2t/BJtGQu9jAu6X3zYoBIlqhBy/KivombMzNQDd6JYRmM4Y+ytkBW47pN
qVvPwKgIlpbqQZs927+Sufb5wLU5bz5MA/zRHVA4PDyew43USQV8RLkaVLMfxPoLocTlALJU2GbV
Cjjonw5lbG/mK5/umNvax1RbaalP2CoE2cNc7IV0jWlczbSYj/7WwcvRKKs1M4eozZclZxR2dDVs
+H6kgyqLWASBQBEF1OOSiZv3nTCqU10pL4UNXNDBFA//ngqMfU8ykIckvwcFWon9W6TJSO0cp4Oh
4YK4XWdKxZLY3DXsQp0TxCSsHbZPDazuKnNcO7Ards0qKFoJTdCJVpeL4IK7DV0ph/ujKbkWk7XS
R+PX9axX67VxLdJNL0zd4L62cXDr+smrFUsJzWjkg20salnJdKZQ9MJk01yZssNnHmvpXM+Vmada
v/py8M+LyV0BglqYxaAQTbZ2wnZdGL55LFC2Es8ZbFZ1o83mZ6BRFX6qg9nmBW/jNXy0LqDB+zPw
ABQUYusHDCdWaImKG4bkL0yEu2wcTHaKPoeM4ceXNwsdtE7Th2tjm0uV8ozcfTz/OSJ/AUUbr27H
D7I5M1S3KJiDZLEMsW9gWtydtkc8GSA8JhpOJS2r9n9KynXfSjAmzlFO+RYtS2w5HQUYtm2ZxwON
AdtHr7qdComNcQDccky0RnjIgU7JRuXAvkUJSqVybPesnKt5h8RzTV/Dn2uuGSTdFUNFQBdUtQRM
QM1cuEW47aRtk46x3FLwIF/Yllw8l1ZHwK76MRJ5rOckAVb1b2aYjoe5SjyLPFIAiuOyUSnyNM34
3N0fU0OmdF1wtTkQX2Z8JUJfXnnE4sPlelhz/fZ0mJrxaMaZlS7wsagfI1YC2GOVT32gnbfgUPIZ
Dz+Olegnub0LWAw0Vti+iWFOgDu11Tj2F0VVnGwj+/kNbF+zunIYMw400t0d+LGHlagsevk0HIod
xKPn94xaA7ZtgIhohoHWS32YNUs13N+RCjAwGcPx5IdvtZ+a+zWgpiBfTGRfXl/WM/cvh7abYp1V
eNtiUQd3dGkkYYieJcB/ttXEnhOxHNOlfgpAPwHV37Xr5BTfvy0naG48gCWzmEL9lDWT259X9W5W
EqhXogVms35Otyk4xD/3t3QXko65TGtvT5xTP0ClJCZ6KvnQ0sRoMQzWtC8wU8E/WsrJXp94BiS+
b6krV2rS3XYI18uSdahMsKBwo6FOTsKrPCRQo5CYhtzol7UDzYCHytRcSFSA8NCKj3tPhXeoqlBr
StbG2uSiJFe9HWGFeacmzmu/ftdJNDDIPqjfQDtqbZdfPjD2eMekfinaqTaa1KToE1LjxDutJEcH
gUDQEfoRABHtqDF+V+RX/3mhVsvJ8rO35z5ZfYRIUQr1TctFvhW3r5LKUo7wTkjDQBGYMMN3CJ02
Gpyjph9U6tXzhlMxc263i5IywcorbbXJ55mxcfUsnqZ0imMKA3E0/rMm1h2PhDLf0YDIoU9OlsYi
eTbWYeC/oKnu1mKBE6CYd7LQfHwJN1jBfoPp+c7wIDWmxsYw09jPahsTH9UyEBje1RSC3BU+gZsF
LMuujrt/NxDq682kIlDqNujBRarBBvy7RS/wXvIZn3j+VanPvfDgu58RmlOWjBI6hiwawBCSgHJ9
xAZeU5BRNAyuVx/iVRU6Uyoy/QfuR+vKuG4FtthSlwHUM+sklWc1ucQQ/gWX4O9FUJ+WP99i7BiR
Y8fLMDngjWLw1oTAZquQ8LmE4mJeioF4NoXszWI0Q/nJZ+8OzAXxavfwyBteLJvRRuvAqMS3k2ga
ZcjRICi/gpQA1oy5G7dZDHY3vW+UQhtBxMithvnvSShb5Bp2aCLpkfgSlW/GzcPrTnCApVWkDIMe
jEEssJ8bnyIv20s0v0fO9tEAatAlgjLkCFWemPaCnfhQQ0+J+oZvhUQW4PalBD8KMbH/qwpyctUX
tuipphy5eW9V1tr6mlVaOQ7roSzPYuqjNM+Zkk37OoCQfe7+utU0k1/N+z+0LzQEVXfy9ZAt8KZq
xqdS2HKv+6xmG2W0AVNWWFTtWDuCPfVQ2G8Gd3tGA2hKIyJ2dRDICT6TBK1InC+il3hpj9kwlmKa
T0x5D9665sByoDoaprkwpiLWI07+QwzThBVu0dYG9KM7bjwwTPpWMZWAZbu+UL9GkE1gSGiangu+
i5y1NfJRGTTB9PoOKSpnXF3yfj5OKpNAXwYLFO+bfvHe3zbDI8ppRrDp94ETD/i47EOOAaW7koJX
u1HBaX7w6ti3QHKi1GxYGSaLcUiGf3joGz3QMwevTzn5dxBX1nsYfVxH8s7IPhY2QVSTegm7EQvG
8Ihdz2sQVfZocA0rAneMj1us05G2qz9k4XlO+1YSoYZd2k7ubdI70E41jlND6tRSPnCU8ptjTw1p
dN8T0LQiitaDvJdYFiGxxYflCl9b+1qh8xqmr3VdNZP1KcSNW3mgvg9pxULaS+QcuZXUBQ0eHb+b
oUb+0wF2lrT7oHOi4Cn7oD9EE2EPtEfjIMTz1RYGArfaSoYuYSnFlVZ2FnlmI9twsl+DNnCbnCGk
tbHC5inIZCKjWEPryMihRfTDgoxFKZMJ9B4+1yNrUB4Dqd/hFsl1fyuVy9b+jPy6CfPH09hdv9mB
spsKWrLqkqcBfekbJlbEfA+Kz96ryKN2BNrFlQ6xbB1F1bs6V81Id9IIVGVdK0ya/d9yss4uOYQH
rYk28LjsuTM/OY7s+dp/yN2KjcJ72EjVieSvhi2fKQoTsMxSSf27YmAFMbhKFStHR+VQjrUffUBP
0YiyLyvCuuEdw0PKImINPnsCT6GT/l2bTtwrlkfkbBULJwzJjLF8zBLkeukie/XSTJyx3Ua3HjOA
xg5+m1gClvihJsRfwmjWE7giUkk1tA2DV/Sf4NQyEFwHJnDEQCc52hM/m2yOfzr2vdT+ziuimA0p
zMsru55jRENd1qFZ9wkRrFv0CCwTKveQMmX10TcbrGsoXSBfEIF12/FTanARGkqB37l/53xTrk2/
o6T/n6N4ueQK09eYNwNdKq9DX/dmx3v/07AaRG2Qzawr75FMyQGjpqjMnKFVoEp9lpf5n1eX4jLK
UM8sQdc/A0LFYRJ7HfJ9gjptCvTrQahkRNi41RZx3w+7e/4d+TeQUOZFT8Ag0EX2y7jd6vPw5dph
BCBhGdgPC/067SBihwmw6HcYs5RtwGtpJ+7wBOIbGEFsk1PKV29c/QoezesBy5+O+GuDb3NzqV3B
poAtGnYL0t866iOvaTy96cVcxjazdeuVipqsvfOcYjVEGpjTTNqCC0c1VqbFkq+4cF6PkocLKgh6
dieCAdOYp09c0R6wx4zVWjgtjAp5fPLI9Dmym/ScE81nwDFwkTVaxmjlpmpPxYq7LnoLLV5qWN0Q
WJknyxKS8+K//YIbscRG33rMEFeCUm8pcjr+uIZr4IqSl8GLu8K70RAr+TSr8vOy4DumELKnyED+
lKRmMr+1lVKKJP6Fcr6vUJMWgYQKrg6AWCbLn8SXwkPMOVOJHYGMgbRgpEisCxJP+YYRFJcRgsCM
ExBO9v+Thb/dzU2epLkAw9SoutNcHF644n7LBJYkvIMIP7Qo5nSRu521vQesKYDo3BTVXA1jMycX
25Eb7AVDd4e+tpBi7FqsIKD7lMADiZ4K6vONxmC8AAVMAXKRhBO3pncrf7fjjHq5AVIjmzFz2icw
pBdyr0HMW/EsCOPjWhEBlIBQ6gYJ6QSH41dJYb4jism2UN1xv/hEBrwA+qKixnU/PjNrB7Ty3Yhm
kAClOcXnEyxg5CTBKvD47tkQMfZobNqoyLrSnWzyGvwQfekG/plofxFGRcXqsvtfyMqi9cG7wH9E
2jTjqOi2xecjHaIerZRjE6fvY/NY7OUZnIWXSf+ibocJ/Mnv/WkN8t+CVkS7ONRQy/82z13bGJk9
0f5GCv1Q3b5nlpSu+YT4KVyFkeZL+yyRrT+nqJtzwSeKcLJeNf/21SYwBVxede71ifWOKWDrHJWO
PdJk5W41J4bs6SBMcCY4JSA43wAnzwlQw0ztBTcjhb2SS5+qz2UayI5iyezormHKUDLwad3fVEYo
UzqsrbxUQ6X8mB4xqzMgTbaQZDC+ZsuEXqkaBmyPoFu/hHxGXqiU00uHkcXMLr2GZD3A0ScX1Zfy
y1mMSJc2WDUaT9c1kFIy5U4OwJ96dx3cZD7eLQeV3775EcU9he5mz9P7SrTcemtJW2woaxCSekM6
AErIJ5zgVqet+86lFTDbw47vxYKZvWGMkgrffST2893bCAObwJ8eZKDWZ+hekISTc/2RmY8VRwwk
Tp5QYiro7FOqBUG/OYgw5SqKDoyEp0kEvIMSARWQZnhBZ0UHRJt/k6vsq3WPLlhzN3iyE7X8pkj3
1w1LKyzPM31VqT7oltWskYJngAbwa44VQmd3V3yKC+s0yPv37JOoRW0gq7tOiHP4OvlLtUrsPbuk
ZMuSb+pBMUCmTeGKFe32J3uylD81gqmOSPi/tzn2pZN2t2Vy0T8bvHZ1LxjPlOjVjNoXFBiLMGiF
PR4dqekoXAFiBIC3E18jRncX314VTYOSyFUs7gOt9lA88waDOICuZAzgF9vLRbgvt97QOAp4a8YO
yfC/wTZuyYg1Sca7K3yfc+Mx2UhX+yjfer+Z85HZSO3p0FQR0OdUTrWhR8p6lDY7uZcrvaYTzcE2
KvaRa2gPbHEUpxURRPZbukFYK3hgkDbw1giY0KFFBeNJiDWJLB5wpdsEkZcwbFZU0PagGr+S83yA
7H2lPyK+vR0prf2UjGNfNo+LmO5zEzwENKIa3XK9MfGT6K8jejgI2jQZzBnmpc4fJQU2mmxV3TOE
vLB2WxInUrWuUvPBC3S8rkQZ7zDGI+WztWesxh7bk4KZPZaHb1xP0+0iyXpyrU5+NUiMttVTcjK5
mPb/Embmsyqm42ZArLdlpmiidyV0PtUKBKmciAJFxZiN95STFFKNwlHnLvxIqrZindTjca3W0MTF
LNuQpHjCxmdxFhQVBtueUm51Id19FMW77IVubd+E6u+Oa6j+YZfWDZrqxnJS+HGMcOjurdsr/zEI
H26Ug8ZiObaVGjtNvv1fitpSZxI8wBGPSU1L6ctFB42IYx6DrKX6vd+Igbv+se2l96+w14xJNnYS
nYiCu6VNpEpGgCWf5qmjM0HJZM+50AaEqMfHHWQWJwlDB/v7v4QhjV6vLqQpe3/ART8Yaik2SLx3
ioZVLek+TMH3oyzpvw/+JHxVsCYKLiZK0pNfLQx7RjHX4jG+PA3FO84ymLiK0yClgLMCzph+IkRt
08J+RVviro8DN/7QGZqawxempuVe62u+bL+J49oOEJIwLe/Yrc6p+2tH9ScPyRs03okj9zRaJB4I
SC3aeXg6VPvuzqVUsRnCOVGZmyrgeRjDGNtZoS5MBgwnXP3niBp0qmxtp8Uxw0mpJ3c/ANLJI4YJ
FPvDNNM0vu+FhtAjUWQhS57a5Sl2htnNB/4uKFIFA4rSxMHjSoQ622/dDD9iiBerQex3kQKp8Id0
jntLuR2qPu6dX2F6T8j3BCjnSUdVHDtaJJBr9hfZ/birsJNLA9ANdY1aw/wtsdvGxyZq3g82+32v
iYoE096Hj2+BuFf3qaWuy1zN71oC/92HixYvbemglhgvPKTH9Q1eBEjFHUq13sHnT3+/yO46tL76
Z3EuOQi97HdpUKMrK//89IJDZ0kXea08hNngyGSyUpCaQkxEFV9UmVRm5X6GSau/HUs9/upqlpta
HmMQQHWhPELAxOSE2XTEN1KRW3C4vIup+7ouElUdgCAhyQ23SYzBnDLAAZP+8fZtVv5laY9B2IY+
3dkTPKAuPi1sS3cBrlKWUknZ595SmzO+p5+wrgH9FBdQ21uiBB4EuHtz+0k9J7gsMNZ+b8CJfwic
7SHqhxXmuSXoi9f3cZhtJWCantcWdNw92MYB9GFlcuVUewCun9pztJORLaJORZjFw2tenOXMREnG
SNztq9zZNgafHlJpev205mGq/Cg2VTqaJ7nQ11ZvhgphzlW+W8exMt3GN5aBJWZEvYHn4+jtRgw+
h1qEeh/SxJadYoDcpj/HRqDN1gbAGOfxGqrkyeUZNtafhx/0D9Y5kCxZm4k3PQwsI7ZAyNh+EePN
ZPejKGc+WpxAqthqmw07X2K+VZhiXo+aXDwyIixI04CB/JDECmCB9IAeKhyOqDJKkpyayJD2L3Hd
XwDR0OB2yoqZlNi+1L/QEzWm3F5szzOdzVvT+SxlLPniZGFg5MH4DL1yCAkYr523rR40l621x6CF
8oMenr1lJ5l4fMT8O7iOWhCeQb2O+w6yw8/JAyoSbkOIX7JJNg4ynZU5lxo6bNhe81AbKuVvGeR5
nQGs42gyF2DcKt/1tiaxPACm62EQ3CdAEQj9kR7BMrVMqp8aWLDRswLrA/Ddb2/uCzQB92yHN41w
uxUcmG77jDyolIhi0HTXToGNfdycjrCn7O2lVwpLfMVzp7Hlezhp+75MKxOM1fBZU1XuQYMpW1hR
p8dgYJy7Y9H96oI2y5j9EtU/VmUQX4prfhoKXUkZ4ci13x8KluLA4NAaGGbAqX2rkokgoAdAL4L9
m/FuZYJqJD2Lp/wguIIlDnB05AxlfsxZufsvT3jK1IvSMiyNeVCPZJyWLg5rpdUz8RY233FvyEaA
yxafNRCM/x6w8JDuAsXsoBF19T5p5/C/rsPqSqQSE5iFkuG1Ni5UG6UOl2HsN9N9kBXrgdpAzFxw
OCtrN7an2PE2bfVJ9iGGBVNyb/HDPakhgX/kv3rdbRJ3S0YihuDhMyiR5FY84GLdSj+pP44BJh3P
ape2Kme2a8a/wOjZJmbqevTG6VH6b888XE7XKKhf6rISzc7Fm812s62aMe+FBlK1ADiwgbeCFr7Y
qr+DA+Si3aGch9SG97uaf/xQb5swuSvVszpZVMvDEXmuVPUZ4al+1mwUOVBSPugr1I/+AvSw2gYD
BFK7o4pnRHzvgLJOB+JJySLQLpNphxtRApviv5PzWQvz6kP2I1s9ABTOSsnt4lb1y4udQVgKe9yr
rulqFoYQn/kFz7S0ARvawhdtSP137rte7MxJ6xxhL6ogyd+exO6qmdChtwlEzMxJpwybJjFEGETc
uAHBMHOoVmxSWxqAB7cGm8IQu1+8mskfkGp6ydwFj1a27EC5Q4Nus7t+kvzksWwGszpZRuCiTDgM
tG7APMpxfn9nHsKzRrAv/TYrcPZpx8olfoIMcg2nDfAIoCiW8ulNrRo2ZS1q4CRuoRdVvtPO3WmY
QqYn+10uJbF5BFEe84+gI+adW1Z9GaU3gsG42SjuCN03z/FM6xfsULcfuwQ0vCEM7Y2304OjemV0
cEGdEcY9twWb6IdoeTfGVjhlf8wEHHbuRN/8uQLq2m563qQNjQqtC/ohHjMVibJtC67vTQRkSTNK
o7patxNiq36+F1ICvY57sWuesUvC8hQFbM0XtYVVATjxajQLX9AP1NBVExb4fVyaHHFLs6lJJ5iF
JciqCUjCpMP95nQJQ3YOr1fYLwUaDD7ApDEklbqmHuMfePzBzBJdc2VYSpvY/iX7jC3JRQyuo17z
FmBrS/irYCMvvKL+V1LyL+53g+wUADzP6r6kbNBAdjt/VFoe676RXdFZ6eA+QPWD9aT48NzF1WwF
1gZ2nRfvqFlQ+rmMSVEJXS+vc45x/Yvwn5V/pXiK7NOe9UUDpeWu2bUXT7KYMGOoMKabZ5J9BWF1
1fCs5iC0zjmzXTQ8y5QmT7RonSxRDTwUd2/WcUjQNfdnOBernVOTVjy02SNK97sAVO2uU3BomcyD
Qp2khStBhz40yhK3ZRjRHdaWSZoJ5q28xNDdMPJVrmEc/lxU0vLytY5ZwRazUJQxBbw8bMrj1j0c
a0hrs3xBEndMx2mEmPWmNav5CwfTmVJIzlEATHKcFdx24Onp9mBw9ykeyqd6V0B20W76wetsGmQC
R2DG7kTA7oV5FTIMGXZfiMk/SO621m9aQogdHll7emHqnO8+jVXCb2Cy7MDLrnYzxz2XWY7kcVBJ
Wq8dxSwk0GnH5UK0d23hxybdb/0U3J7fL2FIl1f38aWSytWH76S9c4QjoNUc0g+Tv7OFt1lDegBj
kASI9LE2CKq1kTkySFTUdc9yPYN+pbGh8I8Yvwhzc8QBkQ+GPSwYV307A2VRqLSMdD3s7C29vnMv
2BqABhStLgZ+wS4b3jimgBZ7nYHPi6bTd+0sHrbakH6HG6GQla7SZHGc41F0sU7Qa+NgtnC56rzA
DydmxdTOJW9AbWwgRxgfe9g2cOc2A30FNDLvjdVkbgWoo5J0ceRN/o5FI2Nn6+2dz9TJ+uG9traX
93BGfOXaUD8V2R/8EH/4h3oBeKJYbduQe0nEWINMXjyHu6ybsNFvMdTD9JV1uQl9iaH19sbqQPSA
vKfvo02WyjdTgVPRp3Amv5MlEOo2KvNNA58LQo0TtHEVIFZmQllBl/roG48g6onjg6Eb2Pk3lLC5
xeHoJRe7xeCaJSk8XCn+USIHdrT+x7a5JbcGhEajDR2vhhcfIu10reTzh7l9NNvbE0haZsFuLOyj
8rY6hApiVTad5r0zeX18XzrkWj/+IR+w9AHwKfiCuwO1ccRu4oUb0UzIPFvOBYyPuznHL86ZpsXh
QB3kiwpp0lQMnkt7URtr140OPWE5V6bl9EEr2R2t/BSSl/zhJf86o2Qrx9VclUQA7EaS62NfiNLN
IJ8eraTlV5u2OmTjWNYmKLXmcIQD+zuaQApfrLqN+EKYaK4W1GUrw62MC7cBS5/vQDeAx1/C578y
OWaBRXVUMxsuVBTbYCv8/eYik0RltWuDodWhX0/LiORgoN2K2euJGteqy9Ui1q/HzQf8sfORMHSI
8WUxNM5bgKtutfKAAlaeTkHzc1nlWO5mr19VVdEvr8jwKkmNnFEXRvtioQpSOD+zkmYaMCnsCKSI
4ucZsu5kDehWTrtPTU5BV3H2dTzHr1xnoF8NV2ouw0kFKlARuPSodcVkkpqyJY2GmvVkk1UO5E8X
bjcq48Ajg+WLUp04GzUvtlAXzClvNAbrJwA8ugEOPiwp08t5RNokpErjBRbEsNcNu/+vc/wB64ji
z9SO8CzzUCef2BSwHOEVRNwwC6/F+iXyDixQSqkByXgY34KO2ngYKb8sZtpEbTBiGDqyBnQxkvnd
10WmG28BBuAabEx23Eq1q86ls40H6A+JP4OASmduBfF4omw6OZA9yB1JN7kN7bQl2tsXn0IofcFq
WsNCKqettcujhXMfHyfIQQPNmDSX+v/FsMY+4H3ZzQzu6K7ZyA7k9LjmwhoyMKj2mBZyZcqH2hZz
81PJYK5Ol03743LG76kd5kMsoGZcK4iyCTCm4+hprh3v4K65MTK6XM++i7rYov1rNpxQb6Jxu847
nhsh51WpwTuW4XByyaZtlLzN66BTTDA1gUoZR8DrDqorZdfFBRYA7ZjL3vuvGMcuyjHWmXuOidz9
SxPili9PUVMJOu7bUSo3+x7fPbQh5eULy2xtP6jItUL2nbHKTTXS6QdBvCQsCJoNZrahjr60VSn1
ujwNbz69lhR4Qhv4oo4D5k9Amd8CBiwMaldRQ+PJieT0+85ShhnW0tfd8DqPQ70V7q+I3HeEYOfF
ZaLlh/4obpOKeFSNjJ62eVBJCYaczmyjlWfiTRk9ODaofb8O+i/+65a92R69LI/R1D6MP7jbw4gP
zu1dED/FJlxug/LsDl9SIc+uUpKbNfsWI61efagVtvUx97uI7P7mb1ddu431Xb+HBMrRCzyETV6G
JuEjtv34Va1zICdWXkbXbfqJ4h7HfNrH0GI+YXT6cnk7gdEoSDPSilEPg0VN/GttLbECDMHwyyhM
A/n4OrTG1tAlc5ktPBGcSg1y2kJkzPBufHcAIaFxACYENM9PkE3ui2JzrXMqcp2n1ZOhRsiGJxRJ
qeTau6X7+v65CeAHRwt4pyFu2WTnxtcHxYht+UCGARFNKy6Diov/LnUtnX5z8scndWIphdDCEFI1
OmzEgVZkw2Sr8IRkbtvd1I9l3p1yCMFn1KavvOSFTScOtLpFp1Obo9n5IYUdYH4JqWaDIaldS8Da
cqqDyEIInvcCNL8o9WV+uma90uTm2MIWTDqQD8xmnHYV+2uMmrfJ95G+VWrlyX+WGg7OI1TZHNBF
r3LUxJ+QwbtuCdqrAujuSSx5I0SUSHSebLPueVQelJ4AsJKQlFQbhEBYxvKrBZjh92+imu+KF5Ni
CSUnyg9SVWCg6IaqADQ7UBFYTP7JY0zirp5+1z1qmD+8mxwiiaynZREztXk9AwDT9NDNcGRXyout
h5Dwa3V3StRAHmaKCvke9R4VSbBDReaTsOsE4vfmVT5jdOnS/tyQiiTzl0pnb6RYYX77lwNs1l3N
3bNAeoFA9wlEo92iOudm1vbBZdY8L8yr6jbfelVIqD4kF+9SH9OayNoRCNTLF7Qjz17qt206gMTC
wnPqTe8Wk4S7BpGNSqdGVqCHAln4eQ+P+vqWWZEn2oguVjrQ0i0+618UsGGA+0Ns0QC2L0mqqSKD
PwZdd5N7qTYxBW6TxPPEdqAbeDS4dQy8Pwum5RC3srtSmJM89l1DgjoeLzFP/adqsm0FCo7Fmu9j
R3eBD3Hcsn/uUudlzSPK9O9vGKbIo7LWJx4Uc+jlCo7cYCRKjghH0IJzUbltg8tGRiZkwtA9VYfE
byY0kA901DrUZ1X/k40e+3G/b3OGEsEq/NApBhuqbOl1UWmOipzeXAPqEGg1tg5kTcsZoLNVaw3C
y53f/mFvCWrZwN6EjIcavOgyx2CwKlxBJpyPYEQgpfoAEZ03oN17H0IXxnOMLgKsgSFVX2DGBbsa
97KHjzpfIaxFRLlWQkzzTsP0Y/Jp2a9bN0PQODsEVnOPCl8cgwLvlFn9lt9aLxgskZvJR/vwIiaz
v3MPexSd4nSeLAPAkjR8x49q5+VktHC5UfIV8BxVO5sgTAHgn6hUQBMDBYg72wxvV/1U26mWyp2g
weYKBsGX+XCEnY5ZVUbmGOqYZF9Ku5fsXhWxMEv9FjPtuzKET+ImT9MkdSnosQtirESLbe1L2oTR
y2dG6JjS+tYrZv5HE7ca+Kxjo8OnXMFN7p/pghoe1qoWcyOMOwPSBfsiJ7ixqNSH4suwce+fJJVH
s6HYMQGMVXPTieDYtxdhdmOkytWb+dS/Q8wp9W81rbVUW8QNHAlgWAtsCg1HIQ0YHZIdc5QukhRj
8sbT2On1pc6Z2IQEj+b77ejObFYXKGXTTWvVx2nLcgHQquwMeVmOpCdtD5G4Pkp5qmRhCVCbtuoE
vk2UsKOkKJlPgTI0sj9gBKKvYSGpksvC11lx+3Y3nqf6/mMWhVYaITbErieeZGvg0THt7Mwbl9NK
vheRW22zj+N/XfGc/gzB5ExAPMWk/9BpRw3UtBZAXQ1KefSxoaLOq+nvJciGYvf1ntF1KJShHnNM
Q5h/tZDgTdfxPNv/fjnVt6o+eMstOfYW4C5fub4AqkHCSxtGMcA8vPpPKu+zm6szPEmPK8UT+51U
yFaaGick7siRgZBjWYjsoPu+C2KxrsjTvu/eRoV+UOo9PO6LTebcvxEAbqz1fAlN4TQqx/HCKYzy
eJfg34jdRbHwMyTp5Un1WK3D3UPOCyiJGDdDlef6o5G/pxvjT7mmfVBFXVEcSxI+ii3tW8vhmg+a
+V0bmxPnNKxetTU9m/04AYCJjpaUFepGVSl/I+Q5G7Ujt1JLw/iHqU6XDYX/o7s7i1acj9YAJn8l
uHgX3IgWfVRGTP6r9evV/CwENSt/njrakY7wZSjzAjm4FN9Dxf+/smsKUiJCtPguAuGrt3Z0ltn9
7Q7dPOFquMLye/3lPaGNmmdxjTGVgroC7e07MRAHAyAT/PX/kIabwJbZw18GK4k9T7q4Tg1NXgeR
xkd3o1j04+keBH3oKZmzfgACgm5nAUNS72CXOJHd0LBLOMTENCkTqtaMcwGwhCntfpNQYdj/LmBC
J9nKCLGGNQ9IigDnR+c8/0LSFS5oanNj4PgV07QHiEAeUWsqq110GQfOHjxZM46Fpk8EQI+kxdN1
RZFtcFS1O49o8bAJFmgrLqAvlSNKyw+oTEhQkG9pfCsTVWukWDS+IkXXSJwYZeybP7ESEdmhbA1n
m7NPKQpCFmbMZ4H6JAg2I/4rsxNDJIUzQtQsQmstKakp6c1d4yWf31bV1I3yDVeUAfnudrW5xQnn
K/LGBcMchVE3XDO8Aq477dEthtDzG3fyZPWRtJXXidoBmRF4M17sEyoSfR/ivBNSt0+pkHx9fKKX
W7uEDdOqJvTbFtd0fID6+frun2VZeL1FlanIlDxgSOwEUgUBjPPp7M7swjF04nyDC3addwF7QHmi
9W1VjN/UxUjUttowvHaG1+cQf21T88sZTTS67yEVbueY3VnXqk0A5IG0Vh7vOohoDg3bDxz+gwHE
FsfYLY7idpst3TrzesVrgsTuS3w5Z1gTQXXdEIb9J+0XmNMeu28Vxi2OPGrs90EjVzE2DTY7KeMa
gIvhaBtPVSx75emz4qmTPOlpJ1LZsuN6SrNqMsQFTeJIBjPZ6He949FCMwju9ljvHICX0vAtzQ1a
S/TxhdONihl4ZUXeKkvGFxt+9FMt4jdDfRwqXmCbUQp/yWggKihkN1Pw3l+GIyJwjKc5g1SWJz5/
VYCj3XIF66Z8y6Hh9UzLZznESoPJ+0zQqBW35tIu0jO77u8/vg9f2PalffR3S6Ko/0OVlvEFLIzK
D6xXB+lfNWp7rRxHiphs8wWJdeF6XBAwDecnpt5WINFLUHIRHSnkS5gDiePGI/to5QMuUkOvliv4
R0refabxtLZA3NGGsdRLf8FzTdzdDL2R1e02/XljmzZxNVjPIwLJzG75k6N+m0/PfdGJyo0suB6R
oqOA/HXkhMgPisvqqdTl0dv7GFJoKQUfzxRoUSrxcfxWMl+aLUtOUyvvU7BwteKRN9w43FdjUjtK
jD5aO18GRsmWKbvV5duVIMAbI02URglB6TSWI5eZVSnyVvnSc5g6xACqdGdFlRP7wCXact/HTkLS
2h6DjNNimq7wy6Ez322v7GbhPqXrzqhQ9GAMFg/qC6OSt3jDBOuPMzDmGx6bGsBjRTqnRJrM//Zf
kmnRkzVKZyyRhnnvOwld49y1JOTM5Fz3cEGDZySzc7yJvVzUBEr2QaCxKexRhCaa11PSaRHEpUHs
bUnaF43cmR/gNPf+0x2HyVapmJxYzNmNHWt42E4NlAZif2QVQZk3TT8M6+syrxIHaXn33baHt0Gk
wXbeb2qBQtZpoiyHePrdShlKUbxoUWdlte/d5xLw+YzaNaHauk7M16GDXgB8x7tVeR1fCseev42d
IOX3tIqai9zSn/4YqXH0t0qHL023ARSpOmgxcvD6CXV3ddDf86iaW6tTcCkPeO+6+ZTkjBfCSF7N
zz9M7bpNbHJMEhNm6gKagqa1cVzK0rZ5a+uu+feisRFywbbKZ3Sxma18dE4wMsUZqf5Gy1qfVpCe
lz/raqhYd5GWpB32GagPNPDuPhKdGbvfgnvElrA1OTUgUM9qlChem8MTFtVp6LByi9oRF85sOjzs
I7xOqjDv7DWUBfCm0zbUXYRWAxtVFe0LfG4hDJoSZEOs+jw3KWgbjlbrxg8VyXoEDXJGjHGUbcFr
3RaIJVaE1C2kiBGl1BVFseM0jKwKH/eek+V86OwZS5XrmjmyeW1P5ZKGJfp3VvHn6ZpvXzAl+Nih
iW5nGLGdchUKAQQY5FDFFOtAHOEB/rIEP580OE5DEr5Bxejtp7+LuDQfkMjY90MA5DPYOmSKxUpu
+UpMtWJ4MZr01tM4PbuZaEAzc87ehl/Z36S8ZgvuPdcZHGilfQpIPE3SFF4Q8oaOF4HX+YHj8ekU
NZ5IO/np0zR6FuQUfV5T6TDfgey5gTuTc0vK0+GA+tgabF/Lcud/JDtz8I14JYYiFkxYJABSv77m
HG9MaWqYaglELsbjNWTUQE3vOoH4j5f4odlJ/ml2+auGg2g4LhtlbQ8ryymFE/nYddZEu0Z7QBLj
hCrzl9Wqe7cIctM2UM9qlUgK3+YXDthpcJm/7CZJvhxBPMSjMiA4U0HyPanxiZAxg4eyZzp3eZCo
TW1gnBD7kz7ccAIeDpwtjqIrcf4e0QVm82b9lrnieRQwK32FGt2Zt5wICMpRksDGAVC2i00K6RBu
WjFHREWWIHSVMdjfxVQ2zEHnDjOyGkZRrOBiGF825n5Gp8nVh121XUcZF1CbmR0mPc6tGbKzGMcE
mCoVFo5GqP7OxFYi9b928/aDoGpywjljJOnWMcb5Oobxt695BPcVioRheHCXJYVhFnwckHZiQd4a
+r10ZXPQBKElRMraBTILThsaXFFEv5DBPm2YboDcxCDbFpa8kVjXHeYXkVS0m0WljbCiryKb/2Dh
cj0qioqtwc9pgxIUMMpIQ+Ky7yOBFQqV3TlA0aDDciIpoPxO5jmGAv0MMk2d1nnpjY4qTCZhnBur
GkEb9LvAX3C5NwaXeSvNraJ2Rjb0ZR3xKmffekOpDu4KKhLeQe+uQ36qXUk/vtFAjF4PQoJTI/WY
fDLPpnU1GxurHegnIstqyW0CardBUNp5eoCzlgOTe8EK6E8q0QOPWLsPAqtVdTsXpvmEXxq87L3z
kMkONiNsPwFhz+pC4WBRtbTOwdfHOs8TVmYXvNS+hGp8dLoxkXLDoVmGgN6maNa02F97PII9A9zY
J9OJxwyHQiR0T9WabYIJRbZ2OUuJxYqX309yET7Q/cJf7uNJNZyuppkCqgKlzJim26hh7ovgMzeO
Dp/Nz02HK7z0Oh2v1yEpUeSNaIQhgSrHtTqLhWdKEgoeS0IEEC/hNV67D59fXHAFJk98BHI86pFi
IPLSuk6Ci513n4akFlALowbD5VHHg+/S7DJ/GXKeg+tcrZ3w9IMRL0F5oWSoEgythDR/P/FAxMAB
EjMi0gR6mQZjtYzz3gzs2cbnPNo0t6Zxb6Yxr2QMBvzV6/aVjS/1mj8iESduE7H+8K4li82XPoo2
h5AWsTPj+GQuAlo821es+bw2O7ZPACkKpJJJ/IxjZ00j14rqvT5I/BK9rdCeCiIZEJrbYBcJJjJL
zbS1bWlRJo3tajZAl9WgwvIaDKknPq4p0Y/nVVstntIpzXXMrEvKEGOZB16vlzOFn0zKLBKkvHcb
51I1hQM/HQddyeL03GoyHwmM9Obu0OnwrvAos5GuB+ZsZb4gteohlGK4cwzetqfxOqXwhI44nilO
snl6xgxXnTStO4GN74kuwJOV4pQEUDWn4U7H8IdSCbivcufYiUl5wrXw5loZFtbxf28DeQ3N8hIu
b5AA0kVpGm3o3YECU97xHWLZ4vxbPnCardStcCPDAO7Gzh4N2tSNVvpPXwSqSeCfc7GDMssnCJHd
89LG24JA4q+ktmu2ILMNHe3vqr/NiQFIUkAGGmg9roKaXCJj1fPWBnbBBJTSnqH+Bj7FMqAOxvSn
SL+A1FMYmI4GgArXMdSF9uzdQ0+DQd29uzjJkv3PO54ICjvN0VItvdjakFI24iGtGX4rc7ket1da
pEk0masmC5bwW+B14Quf4v8YfOr4lGR06YYPQDcVKEmNLvdzjgIfw3Y1KHUlnnsiWzMtXX1H3Kqj
ToyFZrX0gsoNm0jk9CRRmGNAF6ni82JywoeMlee47mOqrceM79vLYusc+lyUyG5IheUEEQogjmgv
JO/N57UUmXEG1+2UBkQauR0n1H7+QmWKMkHnkHT0qEaq5eMF7SUcMXRzUg/0qcoG7+wbEaVi3msq
xQiGd0K1ph0KTlpY56d2I3EnyaUEmvKwNTzQs/1aV2HaaEtr04owX6pH4YStz+3G1m8yfAzux6so
My7wivUeJjILMSm/1p7bkUnvDLcMVlPJIRK/jKPbtxJD4LfBZwxJ98bQgvzsXzJFrk/YYAnwAVgJ
lX9dG+n4mAYui3+s4aOw5zMW4cV5fgJWHIiFi+FBN6HtqthxE8RA4+m0A4HIeQQBYn9H3ueXh4H6
Ljiork3olvZoQchQaWbPD/AMqKm6XmpslmoyAoTXyGO+cO8rvW1eWnMvvyaHJ9qctEsWENtPnG6G
q2RZ66MbrU2RH39obZhZ/DhLlLdGH9ceKbChgrkzwSkdOfIpHdkyMumYsNljdP8kJ6qCZY47kE1l
/32kbmQP9SRdaQ92zDRnXFin2zp5grRoxo3OCtAy3QAB7O+zKeXWTCU1gZsLSD+SWrGjB7GLKANv
QAt7rSgsWcAVrnGN8B1cyezZg+uFn27D1kiLfY+qoFlJGQMh/ZNvqDONOsy+w3nbBQ+8ICa4hj1J
tTe9xwk1o60QacM2ml8C4FX5tSkefdT1/d5ajTQFtLyqbJpewVHDQEYrmDSIdNHwrOOREvO1KEaK
7chF6N2bFtn5Hs36js5/kH10vxV9MkUJ+ouMjAg7vlKtvK327ZZ2phWd/UWtWTV5lpHwF4xwBG+8
MpfHjOxqgh+BazE8SDJR1w/rVikFURVhEUqVYm++K1A/CBi6cyLM+lsOrEE90DQpvpPoPEygNvNH
cYy7vHMYddisXNqXDZo9gcvvx+ERhRov9cVDlUKBD8V3NRklQajTcTfXXWIcXCr8gSW9rCdEYDcQ
coQxUPmQp5/9OnHcrE7nfbxu5mRSbKzuGxRVl3IuuNn/2Gp50VjHFh9wsQxIqkQoQS9F3img1cQt
Au5fsIUpmBg2yYLiF4W0oNSWXmdO8Zgck8OfmqQOdjHgc/CH6zCM19GENfqv8oOy7V3WuPDmmtow
SNX1g4IU62AzIbTPKf7WwUcD1ODWOB/HuskP0hL8FgR64dRQQjttQFaCpghVjf8LeO6SnPzj1BF+
8XIK3RR885g2iUJy+mzjf3DCtClzRii9e3fvlHXfrDHb1H41YpWVa3g9vcATqu9rTRmzcTZ3dJbL
NL2tbSIAZ0zLqkVbCr4TAtkruJp4BxPK95CZthc3ztYJNCqvpvSNgCR2bJTPbwSzspR9NDNKozwv
DEoDwk81/CWqGoOoXv4AXNykkrGyPZlVaIo4cf+XvKEyzHCHfLzrFVzhJy+PjHVzrXcYe5KaFtx7
EUjLvR80NveRV6uPMrpuVAwLeY0kE/rixfn3c6nD5sKLuRreJrFDJi6vL7dP8qyc9z4KiL5OfQ99
WwrEjJG8xJL49cBjbRMkj8u09UVLdkR17PrxLRDby4EOI+76eBn4FyuEDmkRedCzeAY6/A4nE1yL
Sx9wxp5zlFMKyH8tzPAO/m75sTgSw7v4nkn1F/0++jgP4Zr2/bcMPyAXvwREp0KzEVfQkB9ZBdXj
B2sQ3NdLJmEo8w11G2DpDDPhXlhXLJpcrP3zJjO81WG/ezZeqYDk48seirgOylqqRxoHbtoSUMo/
CMSeqptkvfJwvn4Cz++uzfkQKOflz/qOeOqq5ROyQvai9JSHHUOLoePbCUqq6ml5lXAPSVeLlVlN
mH8WZXVoJX/DmSV7Trf/8Y8P9mcZWblD9IgD9pRsI7jwPti+iN/kn6s2GUAxoNjrASLNY+uAxwM0
/eW+9X8P7egBVptSPoqFRd8n7meUX30UmP8aMWzGrnXmNek8W40qd2GC6/pL0mCzw3rIv6gNYMT0
1DgtbM/NkH4VYY4BWmgvdr771e2uRTrwwvPc8aNXxSy88NXpJ9EyPW6ich1W3t3lfVdIv0u3zWXT
cUSVNg8hr9EmInMvEkTijBANagzMOBlnB2CBcr3gB/U7Ig1JKX0PbRRgXX/Ae5jx/5IGSCLfM7Pu
gQJKvy2p5qntPigRI9PgRQDbFxSwpqpeJ3vcqIWQ9+YZopA9t0BQCZzuZrw0KOWLJ2WsuD3VEXaT
JlryUq1fxZ4R+OT6/zZ7oqSunhQP6r1Esquz5rsRW6GBBJfTbj6Di+BOttnTa/O+bUvo8Qn9pKzS
ovcNSheM21b6tSDmsndegkpCGVbA/vMDC6msbTnm0MVFvHrnhpstwwbqf9Lu2HGe4oz+0sJ9j+0G
dWhcsXya+hUDqE7ZETpwQSTwWqCF1vQFBzfp+KtsFVo9hiDIy5sFLuqG0tuETN+3Y13BRktldmHm
WHQEmnt9BZeTynTro9LMs/Xw1t/JIF9aq5S6F2kwJ+bVLjZVHjgh8UMVGceicTz3xnMeLn0D3mo9
qMVONa+DnCBv63BsOyQnqDYHCYC5yEzJi89bSTzy/7DpultcAztnCONO4cqbGKdryBSExhlA/Ddp
H4FicWtV0jqXPi1DV2uirZRfOMdaWnEtZDj4msveYWyRCR7D64zQcmchTGyaECgg469dndna4vda
JK6e9rZ6aarFuSAF0/U8yXLFaA1ZKngDy7qO9bfGvu7+AgBrrFyXUastmaByFZyYv1XRipLyAxmw
xR9QC8qHAu5BV/MbWEC3zdR7hpOoaLYDqkWny2/uO58M9I445503uMbhlb4ioDyD56Vr719F0sCt
3cyEOvbXu8UyhCzfyev+Z8WaAhzRmArf4m5j7bqz4mTCk7YbyJvl/sY4C6xJTYvbQt/jt/eo2IRO
iOJ4jbpqTrbeD6PfhCTubZuo63h6RfOWEfVNu8rFlB4YaVT0u7FpQoZGbzKNEVzvCsF3cyZYzeiS
gc9SyrBtiyj5XccwVv3kg9Y3vn6Cy1Q1aQd+EEwDAJWc9u3la8snPZmnGVvikq6+YrPH7p9SEqjA
86z0dAX1IsIqKXj4h1idgjKPGioENxbD33QA38coVJdCwfPfpWi357lUNY2DAUnfv4EX3PRu7ecE
hRylcXvaLKhtExLs9ugml6WJ3YJHR3sU+U4QlUSUaZysS650Do7s0Q7CU62ibl3Yovyl5OL0OJx8
hvTEkfFG0u01Ehq/WZLY62ENx7W6x0wD228SPymz+DPjZp5/BDJvlJ0ZqXzJxrbFqxq6z+y1/2GG
lEdzzjvVGoXGWTPJISzlEhMev71gvUQnVDVRXfgIRLjnfeWsFgl0fETYwB3KLO/VjNPTu3SDyXoF
RHBIZUcow/OrPwP57WSKhi7O3yjKxJgp9+d0BKjRyWHWhuZNn2BTTMoGEBEa91z1ZBGbOuXxOmbT
MYwDRuqTH3h9btvF2fhafnkQS+esyfPRhjZ00cMOUW3bXLk/BX7EIsNtXe7HDHMzvCh7LLZ2Maxv
5WNfhrdHn1ECHoDoEkiUAZA/aRQkWBF5T+NZ0BDXKoKsEDkGPs4e2lS6+p78eThmn0EdIna9+MJf
iaVcuaV4rpYuGbx6CeTd0RqMhWJKMQD4vbe5Oj9/FKBcGzaQ7tn9FNJyg5i0W2IYW8C/yh0eX0tW
5DN73oL/e3lRU0//kvXLaQxybSl4v1+KuqI1etdq8zKxWZd6nUKL+p8ZlXP5MGhdpG9fTWqw6bUA
O3DEiY/FbjbivcvZASGAa7Hf4b/dU22FSo6RqO6R3FpsXLzkYbP6HaddJ0gO9kdOSC/zVm2ntaJf
eUJo475X8tjKAXaKrIAgICCyIQWd0hX/1+FGYS7xxlKKccNlbeTBPLjvuaJN0eyUX5M74lYa07zr
Xhw1GVmB4GUV6VV/YXTagQXsQlMnJyeDiPbVtfG77QdYHbg26I9r0X/m22IRA3AiKiGMcJ2nwQ2B
b28daPPLQmQ8EjEvXbnBMJn1dtm44FSk60KLg7DjCTqvpB+TErBeo5TOnyc/ZvSW1gZIRxsrHQOG
ouBz7piwTkT2NzCLxdcvR5t7s2ahSvviKSmjzSoaXO9wl3CkqD7zlgS3ByDb0gMBvXiy1XIz8CIN
ZDdI8LuAfNwIEbmX2PymcKoTry1274LjuqMVRDDUtVPVBdKH+Cd7AumzzFqTAla1QlNO72Zw7sxb
vVy6cIdziZDciFt2PIs8D5U8+ySmKEd7AaUrWSE+Db/tBWPuo54wrZ2tJgcHL2lOemo+Jsh6vYLq
8Lz0tCflEMxgw/UaXtIn79FL6kXIBmhp/trClx64KrntTar6TqIHMNWmCqKtLS9+HyiilokJ9Obd
bGo3mdQB5tuH8JT1DKnMwnk0hCdHwfYJnQM9ML4oDBkExGpsaeVWisfApAyIgRuzZImdzDjowGph
0ZACwlfw04BfqKCTUjlK5cBSfcryzYoYaRwGMxA14M4jYuKtbaJ6GkQv5HzNkLuoIddl/2GcNxlf
cLxoDM/QrmoUOx7/18LAltROR3TMElT7XjQ95R0oFOyvpsu0/lTSj3RxkuklZL4FjD9N6g3XIpKs
QYJ/PsM0ilo0o+DEax/au+SBFEVPo+9DI+I926+xXLs6B6hAS274aUzGXtNxhxrzpNNCZGIjB1YY
SKEKpbmlkfAgehVUgT8wlpYycsxjMCaZPpa9XcGKpgekYrPa4MvS1mbCmEi7AikmAgLYl0nIOWkz
ObJ+xe5xk9Bwj8n+GVbtQa2EstyydtS/wp4cWSldqrIFWV/KUl1K7vc9gNsH4IX//RHeQwDLMklk
y7y5w77I86+r2jBIqMG12Uaey7R59aZef0+YI8Bk+PhaJsgZVbrZhxXDe4KrVz+p8UTM1iUerhW+
f7syslBWqXT1bq1WL7iHnBl/qDo/V/mBB0CLHrTMT8ei9rXaNj8hkl2gW7KMjkbANFv4prIBTk2F
wLXw9X9Tf/k7EUcMXmYBE3yCGpeMwB+huUOm6R7znhIYehWpxNqNOT1Hxpvu6o382o88d/xJVSxb
w8oh7a7HmNPf5CZ92hYrACKW0Q1AwN/PJ7xa4AusWKDObzC5zzZRAFTmsWzivabpR7a5N6WgZLp6
Ghh8ZbX63iJpR2SSTcQw2uwWhmPYQA4GIrdZkNU7ZEC4aRXh98h8oc73KqIJs4KnDQMWYJozm/05
CyxfkamyRa0ceC3Z5OV7rLOH/FNyOL9F2Mc6BK/9TKIcsV+qSJJfQAOCxzte6Xl8qtL4rR57L4jA
fvs3renXyFGEcVMPpQtrZNHOviAh8LjMxXnj5wS3TaT9kOKkGs+5BTGtzqaq6JESaZq8eJLEd/oW
ujO82MP65vpwDeT5PuJepPXYRIK4Td5jCUXApmB/SCKCfDLROQ6YGYmmKVTOfLOTcDS3yFrHIwik
Ul7IApPJfN6lS3fGGvRv7VgAK5YmSR/SevIzWYJfdnY8Tf6WorBn8s34UYXUAU1uUjHaG4ULB/sJ
8lVEqjxCox3Cz17uBED/LXAXhWt4e7mpvmfAypTg8BvNKlB3iX8d4Dzk5lV8WQ1UqP0j173kUqtt
qW9VIPhjopC9K54X4x1lZ3krlYGfCRYX1PLUbs4AUvRa42DgRh5jGuxCvel25VjaaB4lnl6ut37q
tiUJUr3drdkacDSHDJz7MQAAVkTDW79rZBu0uMljujtTtDgZjJ0wk6j12N9bqoKHr9Oo0zf0ZibD
ljqwC9Z4S3tAHNZk5wxoGsedSg2BRwR6KpxhhLCQfaZDRa8YRx4E0/ST7v7OA2Vc1hKtrj6XO5A1
CCgkwv7s56zNNy6R5kJnbNCSPCSWoZRmNEXmE/bEhZ7+61yU+FVYgkMnhajyx6iitAEhCYS4PxNn
DR7qzaXRXGhIxczYpWCvCh5MTAs8U8LmmQRCqGzURW8w6o/CvFkbbyfZ8wyiDTgLWC7l3/C+M02i
DhNxCulE4oA+RnhePajJJCoEOkF1pwvOyXRlOMfxG2P6bwdjO7DKgMcB5Q9bItsVadnPYY4TJQJp
yuhWaX43Y+DjT1zXyL4gvxPBFt22H9g7K8aLtva/Rc2abi3p+FO7HZGCZ/HwytKeZYHMRS3S1seT
FyhJ2fYwXqS3HEoLsJBbg4AVP7kA1TkH4zteTws40sjIJPcN8T6gw+6F86tl5fAsYtg7W0lNKUF7
0X3jBZeIocKcu4ZTP+ae3nAEv/hy5tWR57/orMtAyMn7411Ln/QKRLq5Qong5RccID7T6vozcRm4
vs8cFvf3DTinSPWiCpiELaTqhQUtn8KtzXyshaDhRZCT/ywWuRPFG7BmQZd46bDsyjwSQy5uTa5D
Zo6KpmU3X3r1DHkKbM+A1PdG/QYFw4tb6/BRiFt4NXeyYqIfbVQo4rV9h6SqRspgMwpO/m4nTQEE
PMn5TTuxtrXqzCKC4cgFHS13HMCSFolLAV6JnA5nfZLI67ii5Z1apkISpRSlpS7Ybsad78a/U76G
qKOnNbokt9a1Mfeke0UEJJeAqT33VJ3HZZdAKgcTBN0tgiiMWf/9Bv2Xewj6rk3Aj49eDBV6UvJT
PFCrBMsGzmu7uvgC+MSNXdroBE5V+7snKEVUS4jXlK6YTpW8ddQklcU9SIzAFhddxqnYulyBpbF8
E7B61/tqSymzRREzFPgYf0+cnoDZ8eA2auLdX0C4kwSCs1rrVmz+koos+IQggznLI7RKJC4Ng//G
jS+l0AHpyJ/PmeRrK3vJXQDmPcpOahQD6jbe3MXfQJOrjaiUe0NJ7XcgmOviwkpUP8HsXlxz9EUm
HSbgWbkZJdubdNT8bNXzea0GCU7rdWaNvBGJC56N/PgzXFZP1VKUZYs86PVDFhDUqHNT4mKMk2Nk
8XRBgGlVNyw8QrxY99+OkHcjwBdFmtxg0lPKX4N7tT5KIou8MhXj0kmZMM3TYA4x6LXG4zx0GXna
hSmL11Y/U2c0UrBc+hIAIHqwmLh2vLnpzbh57enj3Z0pcYRykFiPKmvyjOw2FOmA882zEAtI3hm/
4osejKSn4dxm6scinyG9wGJ9k+WUzhyueZC9O9zcUs0YGHq8NoQ1hbV+u0JRTBO6Zf/oEfm28NDc
aSdCNoFVWDt7kms2SL6bh82J24PLdFqT0R6VeX4cYIxTmZJo7oAMeEKXTbfFcRwnpyJ60a0ZjXA4
/w2d2x5qA8eF8X3ZxD7HAqrJLZRmSnbWfQ3x4rZvFbT3WXsNJGtql4US/JxiGXwCJmFHhwi19eK2
Vuc0X6PveIGKdLbuUk85RPgt09GkQx6X/l2uKTiMY5anaDGgNVDPzGrHiKuAZI33nO0AJGNGLs+z
oajL1EqJjRjLihozm4aX9ce7ICchEy4YcKDqEg2yK56e+pUX1/rg89DmrllrlAPmsgWj+pm2EQHH
x9HPfWrHfQbG0X/cbQMTEUkJ+XYzRf9cLbi8dWPLk0UWU6ZQK8moUx+KbgYpxI/MsU4Xsqe+9QZR
FGFPljaS/QlhAq/doCujj9id23RF9QIsE3OOgRsTY1BEP1QeTtL9alzu485SoSb3AtqIkoNvrYhY
LTrEq6ricYrQ9REk8PZgSTl/e2czSkxu4IOV8M8MMVv1EMeT4lATmWmI7agH4pmmqttFNw+V7uWO
2niZb0Ef0DF07lOQ12F/Df1XiuP4j4sa2IvB3IgxHdUFQdxEh6hM0eZWjmYHsOBqPoBiVvGa+XeC
DcnCaYMb72bR3QRdNDUsq/E+SsusS3H7WmD9t9+0YroqkYQ3A2zv4SD0tPFF8iuy4iStazR5CFUO
/IfZbtkHNtPGY+5+lDjQq4gg2CdUgj4pRktUruGLicP9IkLg/PtRHVR6jZ1hGFBvB6BL/hjwMkb+
1OkHXgPxwkvuGNGEqzqX1wjatE01TLAGYhhSYJe35delEu4hSO7nseb2kLvfraIwvd4YpNYqkJ/C
wJ83vnnmLsflIQCjcLrBPmYz0A6gITX5vRwY1fcQPCF0pbFooiTQfqeuvMV1O9KRrJyQflmcBu4F
JXez3RUrFKAW/aBJIFv2tgPWWAVUwm8JIsHfZN+riRxImiyRPdSmSYAHNMnKZJJgNy5SKlReqmQn
wWBbulj/AJRKgPV/3QJlbc5nuCXiIAhN7J6/OAVl2DfDLSXlG8rcMIX2NZyTnYxrDo63qWC2sxbv
QLdVflJIx3sa2pEX3Zbln3oORZ7kUb+b4tMBQpzwvCiQM9G4F25lGe4J5XTsRGFqwG0pbeZoQWe/
s3nED+1T2moHcFZMnHZSx3T6fyBsJNBgTNDlyuhFtwAjrX5BDMj4HlKwU8FSdQna/d7NsfvdMVBM
a1SGZorNP2QvtB4+HtODXFQy+Z61ctVMt2iaFwkGSSgba2Vc3R98ztstFfqVwzmi0MfOsRid2mth
jTMgl1y/7oJNScXtkPQXNQpxjESFEReKCCTEgEUmXsCJQFDUeP8piNoQZE/FIudKEh6QpASRJ3kS
UXVkhhn8IOZasB/dVxKH4yFPn8Iqh2bIubmn23ioQmO7xtPkC60vXDTfw+fa0fHgwGKqXOv2rczN
NrWp0sMNO95ZJmflaGOkVmBjXQeFqUW0vjyvEXdnNv7WeFUZv1Ogp7x8TL6rZUPhzRODthCuHT1r
QJR+1WZ1RVCQr7d86h77F6Ao1aclxGVuI1fCclBDAmkMAxjUXGbB1kcewGljQyYDIza33ygOlFJN
Fd0HCQ/GUfUI+aISVog3C3XnBN9T1LNX8QZOCu31FzmDBLv2Nqn++cY2NBWiBIKF0jeaWxMu+B1g
bD5xuySUoHtsFVIY+blR5AuhurvR2crHrIVhY1k2mp64dYCcGIiD//JQb6uFV+MFZf7I7Xp8TYPh
EP2qJ9wmZ3oHc5QBfVS3lxWmqR8RbCxPUuXRvPZAcCG/75sJvFnlujmSzT3ubCyyd77WjzSeQh0/
zC1yNSqxxjqF4DIC7RHauO0f5NmjJ3n5HHS6staFa8EsXPpOV4ErkXMyK/T3fXKnAqXlwdnCE8q/
20VYeKYWnMxUw3hBZ6jlZYjbcZ1jMjzaDU1YOJTnvyb6Wooo1E3TUzQxzHOws3r81lBz7aegqhHz
mWaZerLcTLRyx5RxN0CZaGtCG8cmieJeyDa31gGsYf6qZ6c3Jqxm4NJsYYbCauiafQB9bK5z7SlQ
tGe/R+q4RKMqepY/72QPPbbndeBMqA56vpQlGvOAHR8K9wMa7U1rTBez5cDsQ0JC8e0IE3CcMObk
uLmQyuyIh70pMDcLMS1RZTzz3e8giOq4HUTWuzgO3E4rdMd4CDoOhZj7B0t/ekODY8arOf/VdmF2
CMB2oXQSoPzX7H4pph9kQ/80Lh19Ipz3f5zXR3bMEH26TnZZ+6qKmueS1o55/q4BC8q60ECVnfCA
OxE2Nbqfzdim0h1vv7zZ8yPprMUwqXoMeRU4eVP2uCh0prrtYJ43MjmR4IWFUZKDLQeLK/y2t45O
8/K4hHClR0l/X2ZBS6vrfsX+C12TXaJn7RXPJYIBB5EEX6YtS2WemIbE2ZfFtRnpHa9SgEKP2jmx
Mvk1EEw+bIuEonsji6ONm6zG6S0j+nO504UequysJyHYBA3eSJXj0nvAsSJqLV62bMFCLPfV7CQu
R6xnC6YNlEvOoeSVsJjRQwTYCMy6UQ0GuLyvusjRE4mrA+Qrgvb0P4oBneJ/cuo8T27cyfLxsbtU
OvblJbchmIUeIXkOdXeIdsZhC4Z/J4Hfqj1aqGffDwsWdpGI1cQAvCIBHcuZ4pVXKnLE/h5MCZ9w
eKnN6zGlHY/eZm9Py5lHTouA0eAei++0dWg+gI8vHH3txdM34oHT2IZElhoYAjTOXtM4aNIin/WA
c6cWH97CfGz8MtMuTM0QclX9TCZ+wZHqFc7jAwIdmHETxQR+iF98d09f8iy0+kFQDjnZwjQ+/PRy
vjKhzkgj95sY0emByYz+tuItqRwCzov1g+SrycjtTmynIoMKRwHy7Q1btkNCi1aNR3sYJhPmEnmk
GYwQ2ke8cJCkQdTZBxLne+wt6bG197jo/6e2SO+y6tHQ0P2SMNskqwQRS58mlNtShP5lhRpInuDy
4hLutSxAXB0wg9uig25x3e6HYtdN1unAURKSGhZiyF/oBr6pA22V6ONrem7s9wZG6cUigKRpGRTL
ViuZvH8aaE1UD25fQvp2EZ22LBG8XbVfAbdmkZb7LZ/4kEuuq3jkdZ8HROVVeRXDe8C8ZcT1fPJc
YegQot9KZ/xR3W4TOkkUgkuuKuxyvDmF/U7wRO/ukDPGS8ajYlBABHm31hT0OUfWpV3ywYeqM3cU
Wnic4eOMkrefeAl9W1TkRCIuvZ3Kn3+tV7KNk1fOCYSxyUhX+KlWIVtBTm77b6t70UtQpla2XsdT
IpoythFYY4dmi4pEy0jVqQf4Xy8yQFgBZ7VenqVb6H4EyuRGSMK6Zm72ML5rRkC4BSmjgFFGzbNo
+J/xnZD6BJqXVr8ZXE+yt6Le5BTxGrh+gnC2bCUbTLReBG47lUZWoYmo5RmqRqj7eRAqB4LVYOqP
K+bAGslgHNodpe8dK+SMmTTyisJMdaEGvyk/Uk1VOjGflP2cs5JdRAnm7yfa4rabndpnMl8BZFoG
7RLdqRkNjJ4BMhJXIFT0bKj8GzFWrRmbc+UGfyeDBhpGvBIQeFxOklOw5Ihcga5Yi9qeu2wTpa32
lIMwJw9C8WJgxdVsKOs26fiWTEnqifHVicmK+GPT62rmNmxukPtqjzYGQ5dzWHaGRHqeWi1PlZH/
1h2w2UI/kcX5FShU39KN9ql6ImK5b6vC8RYdYa10UkAQQr4CUBrvBK2VQ5FsnM4xITeL8h/EEzxn
w7dGpg0Y23gKO+SHngQue5pn0li1yRwqb0vramPvk2xsvMgjTRdcmrLXIFFuuTPU2yANlVEr7tZV
q6nqvnEJDQ5BjnRj36TD50mvEzqmzWpWX8rieWKOcHCUAfNYGtS0j6mhdezVp1LHUI4GVDE64I6u
TXEHoxXweCOqTVQsNOJHP379Whu82ore2F7hTQ9U/vSSlL9f+tiCSeQHWngdlnOnMeimWNuxFETM
3mu0P7qWU92VRieHWlou+lERDuqPyqmmR6goeIzlt3RiyWGQPfre6ztOGU8kR0eW9vqSO/R8n0M7
wwchjRtIYVg4ah+opyEzjeiNto1Hio90aCrpI89M9SyCfLQyt7kuMgWvYOKyeZtp397Hz7+Ejj2i
Ho0/JbZZhdUoH8Srw53tpPGMCnX5L99TMQXfuu2rOY+SpcwAVPZ8YHO9r4oXE2Kio0Yv0FyP/q4D
+c8/oYKcUjk9aDAEDTDgNH4q9lLkT+u+ML/oDW4jEICrwZYiY+2W0Nysa2lZOJtNd/pHwEFj8uTJ
NAxCGyx1HqoXZ6POy4qKAPLNxnw96AH9cu0Yzf6Bk/XJLCN6S6aDOOkWXkxWE6bNk6Oy3Rt4yygM
shSuNUKQ/tmSk7zIKRMPjFUJUzE4qBhsbu6UEVOs5wc2IfQ2X+S0sIPR9uEZY1sQsMkfHFXUQLq8
axY5+7dYGGXmUb/+Gw/eQfuQLf4q70OVCIrgO32zR5fP2vYmW/s2kmNjwugRmQVzAz5yGEKU96jW
seDHn8dLdZ1OVfxYrUsDVNHT7ujWy/GIL1+dIzlXb47r+nQshT4PUxQKsNAVEy9TjXIbgrEmHtNc
S57sipf0/LJ2eUX8kM0O5r0utiYvYhL2NRXKqHyrTdb8dfkj7xE3aAmaRe1Rx+a5jup8UOp/1km8
7Ep5dT6JzW1+c5VfdSArOrVBk66KsyrPuxcRi2gEBfppl9p6uZSSaBpRxPy9ck75JO82ZH7xybXt
qD9QndkSl5mthrGWUr/hDMOm2bTNp5fG4g2WyyapzF7Yzq+gedUBOhVC6ncVcCPOAkYvOnU0iIFS
11QCPP2VUAvmtx5QJO15jDP6VBidtTw23Xr8XGMqugikQK9rembCPOgmkHKTVVnfy0YlLOYpmD6G
y3HPTn10/tUAXCU66uiheaKBo6FYWL5s6WZGQ1SEMtRjWoHhJXq0uFLGr881cZE6ysqihSdYMtXA
1y2GKmeSJA+0icSeVATxHjtpdHS0H5k+GCyABqgnoXEf5je/MAhDp3Ogw2odJLqnz3nfwrOXD8oS
UkuCk2sXziY2aPxQKUfmS+wWjfFjG85Qa1MukedfHPE/nZWDXWqSiB7CXOGaNz3798WBVXdglDl0
6NdPUCHdDv+jHjr54KB3dW+v23bXubUpHukICgRsqq61suDR8pJH8x60io6ovB8h8d/D6Lm1jcB6
KDd11atJyXKiKnIr1OCpdjWVUh/Q9p8CW6N7DBPKjEbsxmUDLg/SQTQE/6zYlFmtiuZYU6+K2xrA
Y83iHuqT0V8bzO80HL8Gb7dtaoLQ8F6A1QoeHFJcUQPkM+8JQOF185nlgbW/ueYZWHcZ+ib5ATbm
q9h/xfhWpgJTjbVusOlwOTH0ZF+9S8wGozmdghWIlszdXN7fhiD7ymRso7r/5WsDMWgW/cs2qZhQ
a9LyCKABdB6Hln3LOG3rGDlCTp4sfA4QOl2DTgHWLomATpYsWvGt6FRvFBVvTdaivADAJUeuS6BF
A5iJ+Wyw+TfGDnuKtM/y9SWnSbxURiCrMobAJlHpWdblb1G075NZoOb+2tr1TiMqc2PrUt3tavM2
X9jUg61VeyFT41k4maC7o53pnu9cYfF9SJBnYxOMAuAsJpHrdZqc1qLmOoGERIsz+QdCFUGYMGEU
YsQf0FgRRVfEP8jQFsRS7rUcKlvHgGuDTyxJjhhzYTFgJobkwDV7vkZq4m5058O2mIy/NQMTKfO/
DJqNhJGyN3VRo2s18sKMXb0sEqhuSKmlOvq0g1Td2eW75ihA5SUbdYX95+i3QDdvNkez+9YBzv/K
27zPhc9x9UFVHV29WeIXqV52TeaGvjAk6sgVf1WpMdUZ/jXoQN3dH9utUDSFw6VeM+WoAoXHI2ZU
0APZJHhoR+HwCXTXtPx4Rc24fZxDTAW86Oer2fzzJ58YqQh2HQwORzN25pHJL5j6Gj+ewkYN4zsM
rId0igmlsdRl08bo2nW9KBm1MJPNcCi+1FamTWok85n4VGD+zYHNWX/NOERlemrC9LN4RYHrwkAG
CgNGC7FxVYj5HJ5sCv48p5gHOr8DwLnqjGJdKkArmumuU10JYQDeEK36xQJ1NFB+IO+/OEmtiwaC
R8xrj+3vg75C2Ccb9GzU73h6ocZTyzwiRiLOGbf7QZnpH07YTJgC3lcTstq5hPCp5TQq3xyevbqY
YvcJSCcHgjmE+AIkiKNOW3eR4ssJxaqM1M5FPVlHg+mlhWXPZWldv8WGqGPuPtzR6qnvF5MPd+lQ
1e7ixAVqWa6XtDfVRCKnq2GjfnFiZ1WCmHT7rwn/jSVM/jl7Zx1KBReqsteYahv8xXXBjX+WWz8M
mVG/D8D3FEIorh4m2jNXppPpqL2Hkd/CXBc2AzWLU1yRA+rvdRLHViVs0GPN3lrqS+pPjoaZaHms
zt+9Q8UjzbSY3DyvAevzxNmaBrPK9jIy8HUD2P9XtLguxwOPXAdbMqDK45wSxmbSsZlRB77lVsB4
lQA9fIpXD3dJZqrR25AaarmooZ2bPc49RsTEdYbUsyyChwTd2yWwBoq/HA27iwpjD1xXqbFgQ61Y
8ZYo7IVSd+T0/1B4ap3T5QA0KMv7907zdWS5f6ACtPRnjQwRIJqPdYQGdiS+UbwKx9KU8kLnpgrb
vCcMSge37uS3hfO23HtS6sAvhDVqM9yBY0k6jvlRwim74TSWCBmazy/glZupivYOP4OMuLz1nC0z
5Qi2dKBZ3nPeStrF2zcs9w3z88KdRCUvKwaMkYPU0Xy7hnBR8Q8UHZAuU8eyvyLdM/2JA+Li6BCR
yb800KwJbR8b+uWfMT/mjXXTES1akjCE1eh8g68m3lSIeBTt5Q41JBwYbiKHWtQr/NTHjooi+FRg
GoB9EiEpbFIXaW3BLG/wvd/BrwJk2hrsrffL8XQIRH2Fyjxt9RURgwRAiJxx2AW3FrK6si4b3ekl
QO+6brklyFuyYnwx+LZESF2U7qTA6UBGmWhI6IoQ8FAr4f/Iot61qLz+AKPeWchstmPf3WwGfWXP
lb5kdEfNAEqSI83acQ+nYog/7mDqZtXMHXMvI4FrORu+EgM1naOfoQdpbL9WZV5xFXQpINYatWqw
0uYoEoYJj3OjO/V6ysm2wwVDMlXETNJ5tRjOcTX0gV5sTT6z5qhmflCR46w90T9CbvxvDidW+L0m
CqRbV3Rj3243gVxm2hPQ4aZ0MaFo7S0aMlPRCjyeJZ/2w0L33aYeKD4yDyRkzn68uyODmXleZFY3
THcKFXZoIs1OwSZZAGgp0rgNygU+NWRM+qwCOi3a/K/SNsxFZCVZ9xYPvD6Nm6s7oONRF3KAcjN2
NCC7tHtijy8UqKBacLtEHpseJGXjb2ruoWTUK3CwDuCkDwLfs0XRgufsBiLxZ/8qM6Qbd0mRCSlr
Eddzban5fKR3kuDoDdAvh8j7n71Qk0It4RW/VSvySQZmOuy0d5Q6DI5K8/gxsECyJzymd1QBtGnj
Kr919W2PDyhcHRI0alLJaUPJpciSs2IpyM3f5dEQ5ch+/1D/HNQUACoiX34/hL4logRtz+i8l98L
fmXJM1BoNkqxcrTv3erL0IA1LBhB+8Py4I9QP2++GRA5WvVc9e23ZRC+opxCGG7WDxWcBgfcvM9G
0B3t9AGQbsdHRTsaIS5YyHmIi7byAvitkbd2b0zpSkpB6dbeD1UIueExT4B35HkvxLIwNbvFSnq5
mPepAR4TYLRSyK8ydVyEOS1XUnRXBJyxYmx0IvJAvq5xEbYLPTnslJz46UmVYF3ocpUp2PGAgtMk
kM/zRPtbCQky0zCiZVRk/IQZ1pQsgHu+NJ5qh0MMczPj8/upTtjjpVA67iw/M0R8GuoeO0NBPDay
br95EPb82MjAsbmQkqRjmM7kLtnYprjLP2rQA5QzKXUlSVItOT3Z5JfC3gmk1oscO8Qaa2qUI+bO
9GZGJ87Pa6MAGWJjL2JeJCJygq4tBpoBVIxFCkKVhB8ZBYG8Ms38axgh9JirVD2tbiNKqKcjKRip
9IhRuAiLzVXiUqcXSvXOJsdTcT+IBCVg98PoF4a0gmBDs8o5J3lDkwgMUJkV4u31W/FQbkav25M+
EryR+L7iCyNqrWP5805Xs/c8zDTjM4ca2eF6MSJgIFgypTeTrev1RVt4TyViozONFZcc0col9vBz
wgKlnft77/A7NbhTE5gU6lm0EdEiiBpq87a/7+beZ3HGhcP5IgP4A2uMDv3UHq/VMWMGQ9w7v0vw
TG7IM7qkp8+n1RUBShVBJeOjpZKb0ODG95Ja0UeRm1ont0YHa3IamOORihJisxg2qmaNyd/OpYB1
l0rtXTJkdeOJRafaXk8lI49IR1m+aQ5v+PkuLa+ZKiSB4RIb0c07EUPAT8vFVHoSL01cCtqbrggt
yl14HZ7MfdOTVjBRLJXsIC/ikV6bCPyoMgpaIWUWFpn4PS70QsOUprxzA9EreiAID2HSC5ccPzy9
4JcquizYxakQHdzD1hF4lpf80oyCU403WQ9zvz4YwpK+ruy7khErht2DpvfRbmeL6HmtNwwVZcwL
xiqIb1OGcI1QVP3iooP9NVUX+sVPk3khSAvDxNV6Hiks0rXQWgJX8jRct+pQXdPFxcWnj4HGQYQY
PEAW6ELlTQnnj66p6m1WZE9T9M0C/GgpST3YmAFDU6OI5XI/ZBoonVk24/+9iIQK7EcxrzgQsZrZ
INfsJtUbqGaEQHEDTeokKqMFldx7V03c/96fv9IvpabjRXVY5e7qMpmb3hdPi0sS4lP6DP2pQLQM
57xDvh5CUZqkA6VWZvwlGUwDOwHXG0zPj/+bh31QrN8oJV+Jy6vpGtWpWTV7hAM8Y63umP8xir7a
3wYfspTkiNaEsaEKDdsY/luGhY9CWaPN2lD3uSd1wGtqlpDEbkBjEcbp+eioiAAARsu5vJFlDBVl
E7mx2ZECU6xE7gwY3xcmqNu+qZLaSYF4ZnXKWtPu1wHow9Jy28wfrI8Cai9GYk4Wz6g+eW+4IIU3
s5lCVvWhELMF9m/1Z2Y8fuVuyfc4p/umdLN9cwpSo3AKDg5hrXWntuXiLQbU3AI/p4Jj2/YwH/i9
PUSlySjHrMMDJk0aiXi/4UwNlySPc4fZlToQC0efbba5u50NVd8GyeiKvrKHVuglJkX25Ko3qAyP
RcMJ5t2lItZkAMyNkKvCnJ/LX9USB96zhvP2OUJLd2rQ1YjufCI5lKNsSR8+G3qKGllD+xd3CUk8
9Rb1cduy/l4cwmXHF4o/QvcGtj4AQ9LHjKp2MDv/5oV2FHU1GmX/3mhgz+BCHSVe9o2mP68FB9Zg
9l8F5kumB456z6e25jp7v4CIrK8bwJyTskkXpDq4T22zzCbjymny5B7BvNi/BkEM4kUnqNKbfCGM
XNB4RIbgcjpkrB1YjlCd23bDU4uHrnP86tjNRSb+Rrus3k5j3YuZKlyIzPJlWwQDyVSycXamZ1lm
nkZMCXMfOGZfdwRxjL5/l6ybvc4bBiRwNqbl0xsrl/rt7mC3XQkEIYZbfl8SQpf9KFUwMXtp727G
/oi5gr8+SOPpW3mYCLHQQ9aQ7M9Yaovrodz28vJUb6bnAFbGb//8TGwkpO8CTth8kbIkLsSUlwQf
CA3RiNnfOpfKfbCnDEAIXyUlyMz/rWBRxeT99+i8wVCIDfxL7+kf49W8OyFJVnLonwLZKXVO74fo
XwdYHCc0icZ9CMfD9zaeJpFF8/47m/+TiFrjrMx6I1pM8Y+RbEcWiqK+n5lzgaoOJzfJIUO4vcsD
CYVipZ5dnkIdAHLGlDMPOd+YAlfbwni2Tr2YAZMVMWF3z49649VhmEzdzublzvemFxCxu96FusdR
dfjTmrwQEnc5tM+G834eX+fIdhlKJ/9g5ibSZF6TepMawfUAv31WGVOkO0/pieADNvI1OEnybo4q
LN7NczdL9dUdUClTH/4Nb5XSOJw+Q1yC3svl8WzuBkz6p0tpDUXLQT5KDEqLLxUGKtpjDYRlsSM5
lhNo3cQV9HkyhQ/WNojrgj4ADhEwOOPTREDhdABTO0ltDzEaWP6IXR7DHCXXB3EzwSbgBQRaTAlh
/I7hJc/KmM5SZoxH5pMNDc2LL2bCk+Dz54dggJ2JmLMjk+xIDpQ1drjZI9+DDT3k+nTacf+Mt6rw
aSMBRC0nV1Z3hI7PWOYtByw0vuQbfk6JAsF2POSSWsRMjd0kGSNY58yittiXfSHphXFlxE9qwe3y
+WVVhi53BEEFvnpHB/UWC+TWK/bmZE5ZvNNMaAxmWSwFa0vlW4xOlCanglNnA2O2beyHEx7sdP8v
aJ5fJciPr8JkzqCJ8DCzMU8ArPhy8zLzTnTt9P+2Udz9UqVOy0JcVxTO6/rM/Aa/10XMbDRHZPbD
R+mcxo3b9PPK1Bkit3//kz8SiZPUdUWvWlxknGwepeiGExIprsj0zYneAZVPeprryE3VIodXnfpp
I9SONAafptcuQuc/3FtimiagNEkRUJ1Nal99X9BEWc0OfNvksRRmWlWPJYk74DJU3kemovBBdgY2
z3LGxDLHupzGjq/ifLpCS609aOwALWxGKsYkCLjWy4cscMwPM5dK//w2RH4ygUPkWwuaFu3rdiFA
bDRQwGxcBpL8Ez4t2suq/LgCnegYkq75iBqnvFWX0LrPUMuJJ45F8sMxHUzfpS3vAcWHnxaEWy+D
VVfKD1AVVbvhFPEo1Ib2Q+Klle+fHVT/LGrZ4Yhzc161Gg9KY3W7bzc2tesGNwdy8v25M/RtlVZw
kWg+xTlmk++d/16rXaUOE73Aev51jVUJZ0Ol3b/kugVmUVJdQfhawLs+lLsLttmJm44t3Egju9LJ
nnqZyF5lsjb6GySMjf9xNhIImLZqsarzrTuDZWMf6QplZYKmm68gxS30AOEaMIGbiESVCbGTZIbN
o6do3B3+mwCO5E7+nOktCp/Rjz5SBuMAPu1pzMuC0+rO69HI+fiGzduCpLPU7Iw5WI7TnRr61XfS
QybKdinIXKYskXI1UxOrx+O1+hJIsStbwNu/I5DD5OIR7ojlkqCqmgmJ3LFcIAB+WD8E8+BJaVVb
U45xZaqvy4O/mzbE0Vm6eBj+++zuvYkE15xZfIUfsbN/S/n4PkZvjijuq7WGxTlUtD4f6Rruaa1N
JCmLtzP4+OnVYI8sLn0qOPQQGtnvcEZ0BiOXeUr1rFlzKlwg2qcz91xUZRx8PaZ0XdUl24RqgP1n
rvFkoTenQltXPzHcjl9IvBt8N392URYUb2G79AM4E4XPBBQvQFfbrBAKlP/Nq5SL7Rj48i/Nwet/
pFr08/i13UnqBLG4C9DBJANv7GIhwNp0Ai6lNY0+VP4Y9+kawnQ8PixldgwC9xAUXOfgM952bKA4
szKHwsCQbdEPxcWhoamQgM+zYnQZmFVkMej2JkG9TfKx3pEjWPZe7uSFIzMamDjMxichPa0gpnC4
OAWJ8sKHSv9amcu7UWspn2LkMBfauJG2pSms38QpaK2F69mqtLqpR6as0AbnYKsxcDbKM6f+ksfp
OEVAZYUbEHUM1TE63tuRtlQ2mgUjWPd5Su8ryc4VF5Qz2ZD+Cw6MD+P02cadrOkp6c4f1cUbhFiC
YiJiKknT/Qd0h4tbKy8bLEH651uGvp3QKruS62HPzfrYO9RzL46Ukppc61FtHi/TNqX/KbzRU1Fg
CmgM+EVI8yzltbEarCqlvveu33shCTxn0zk8F3HQkOPUVwBKT1sQ13SpNYNlpmR8bHdvfAeSHFhV
SJ2cxlKm8LnYljXclxuBwJZbBVb2dnBhE48xcakVByYpvdRKgF5gh4k1BF0pmpeTGYyvzEFkP5AI
vqjGavg4FJHm0QtQaTlfdCs9PNv/DxtVKINa8RrCi9kvzy4yN/ZmyaU3LSt1d3XF9pJ/yKpa7pMV
cr43vUu/FpdkIgI5q+/+d/tOZ1YpvGwCOptFeh8yisK2uImnm/De4rm/89K0MRl618ff9am/h7xN
myeVzFNRL0q/EBEWwDgrWL9xjATPE/rdoWPqI27/ir39ty1whv5DcqSfRcOGWuEFGnCCWbJ10DfC
yN2r2eZqJtA2+oEmRC6APH32uKIGPzw0WpuoJOEk+DNVBT0jt9l8ZEgCDn8ZnM24ni04J90MWRdM
T3H7N4+ZUIVsTFBz+jJBXn7F0X3j2Niq8MzT2K7kyhmy0+OUNvY6CrNZ1IXQL/U0il4n7KPYdHT7
DaXl+uQGxxdAqxiVlgN6+u+Iw+uoE4MjO8krWfLhW5mTz0SISjbNifpgm79tC/KOGweZxp357kb6
i97X92u+cYx9luFtdIVA+QggtS7O537iJCqTgslUxjVOYzgMT6+Q/E1g48U8wObGbXux4OHYbtmr
wSyAiHnX/OVUzlJ/AZrl+1MXAEwu0/iInPeFHZiF22/P6nDxnf9/Ung9qZtw4QalaQY0p29bEqlW
Mm6tL5/zw4hnEZ0cCYM6gDwIglqsXn5VonwRqrIogJcUdooJ+IaFZOZ+Du8/uEF8VnrisnXCuO29
VQOz7EW/C0NxLzyYr+BQCkcKaKMQ7M/KOgODQD0SX4tgpHekYtAtZxAwdIxZDyNzhPrYR/VF92Gt
GoPTOFAs/LQLZIWazbnfxrNUUFIYTU8WmPr+Xoz0DHnZbN1VIoniZ3uM5nEfJvBDU5O0OGArAlIf
R9FO/wm4vFDRzI5aS9J6efn4mJv/0bRVqKRNs8HusWBaF64rnADL7/Q7n21sFBBsOSxoOgn4WCLT
kgjhOrGdhYUan/ugcxUlitqb5xoHDHsrf8ra9V22s2SH/0vKF8klTxjaiD1OzWZJ+RuCraNuudv3
IRS4a+W/spjDZiDk1H9d8E0V6phYxLXcBx2k/5Asntbv47rbYL7LwCVD7x2X3ZXX/AmFpad3/HUD
wwaZwvQHINW3JM3sUKDk8qoA+19feqOGH60Se1rIGFikoGh4LPFLkRD891mFjgCeV9lMbUQY2M1w
xghI2uiVeMDJcSv8STHV6bGFo3B+gmzXKL2ipcU2dDaaMswvwdoTtot35SVvJadclzVpoBBgi5aK
gpkrX8EKSWjOgsqXFRCMn9l/WDbeaV3ydn6PbGIju12CROAvwtVz1gYx0n3NuBKZRU+k/j6omxs7
0U7WGbrPZ+HxBnyASB/vBCzofRzJ33TuRslM91oXOvk2KsFC7kpAbJI51QjlZCwnUNHBiaK9E3e7
ecSFEyrrkDiRo3ibqwngq52nrt6pAs0Cq8ou8TWLEkOG7a06oAZRr63Zyz+Nbdfxg3VDfvREseSv
2R7yOulVJjM6T8sfm3cIQxemtAcs5w8QvLyi4ZeP0ZL7E0L6dK6nvfk0LjlbecwpELo256xcHe/Z
07ZF6ahdBfT+pCjEsW1odUxOisYOv5b01wAHg0eTzBwCWHzb2HOFkRIYbCAGG+xRcWqVV/9FZ/CM
O6+qgYK+Bai+x9ZE0LtkCmveDUBULiC7Gz0gyqaYkBVs3xriQFFUIwp6wHH/0aZchUraYiC+OmrR
uqM9R39613GVnIm0yPfrj9da8n5uAzGxffn9nEmROY0kKfk6ejIbmJxT6i7rkeZ/4fZuzQA3oiVN
zD0M34tAQ5ld3JBX3/BW0zvNTvvgO8+D8pQyH9KzCIDFbTwB98vv67NO5az4wtCzIQSlEgIPfB+R
ICLwObvJ1XRXZW5dSNPgVxbFYasbt2Ao4Ol8v3KB71WS0e6JKiq5OqZu47QLRY2v40qUNryxk0va
b1YgnzHhYPf7yqAbv27rWLggXrc1BDoPTE1Crf5NPf6Q3BQnbXwrGONz3ZupttvJGxlFHs0mIouA
a0RUFqloQSM8C5bINLXZUmF/4jJHXx7jQtiQ7NN72uILxPJGVM0PxqIle8engHGLcjjWfvgmhamm
SMjhnVVvhP6NjZ6SRGCeM0w7TpXu8ois3en2pDUltjDtTeS2hSalfZlNiDcsvit6jOrHGisGXwL9
8kB/nW/M/QyjS6Rzvl5HX2VoxWKl4/gdTaPayKRe1C0kLgedvwuOX4hqXq40SHCX2P93uDBSZL+m
L/wtf9G4wYOLOrdIPxeHupgDuOrTScdcqmo4AVYPUWAB6W/9nKG+auQYrJyBRFIkENxkfbC+LB4P
Rxz58ihA+7Q/UNm/ehosJxEm/BZFR3PJ92ICCqanDgFKAblAD51vQTEkMzaVu788Tf5D2jB33N/Z
4v1boG8KxUw+sGlHmFNjwPaZXPnk7cHHhTYLyeEJJo3WCQcBu1iDNaxMaZUytGFo/6uay28CVQ+q
wuxlMbWLWmGNXQVC2ihona30TprLvoU4SSlHRbk6+0K+/ewmf3lYXzMkNjfPI1Z58g6iaBQsyWbp
tJW9UQapdovDaIML4C1SkehX2JObMI86nRZmEfyuiCoja7MaSi5C95L58NTLkKsrpjGioaSgVYQn
K3I/TGM+qzZuT+u6wVtWqrO/8e6/igwLIDDsJxbegUjlAww5ilZ1FPCHiBN+2dGDKGjCJPrIvb80
jilQ7yeGWL4SVVbUF0L7p6uA/amwrySyNR11tHMr7Vi6YBT8/5ueX6b98/fH6yqhZo+X1OuTpPUO
TN5YgDtouDW5NHJtgkGDAuUMprP65cWFfWTp+0bhSEVNg6l41vkz6+J4bkA+kMwIg4lVbGZbeFah
fkR7MyjntKMcbpltt3VkKUu11o2ZAkK6KwXLOr55WO2YF9pLvsUw3TtQJO8SwnPQ1zGUliNJd6dG
OTxfPnvxgV8JZww1ADG4ulWpwyFyBbV7mzhMVrV3Oq5Pw+cngT1Bi/dmk0l2sBti152OQPQwbCrl
Cae4QXWjEU+49ShRCWAHeVMG2zEY8Vfoay5IEIJiF3BScl+V3I4WVbz5ljJgDA59FLb2YwnrSUAp
f19TzKuKWsLsidmCsAeQ561ZfxmFErb1wF3DBa7kvq4hqJbLv6iZOh/wiTUE2zFIlXiOywjWcQS9
wNNIKMWKfAFVsAkaXShV5K8w46CeEaMxz2f1ZzUALgNjUXk0v1J0XD5zx9wQZQOwZ/4Tibsbfi5U
DbcStyjtGC2g4oLevQXnGZjPZ7qW1nUJ1gE789CPO0fOt6aKm4/BIurVmtgF248HoItbANX+4y5f
D0MaGHZou3jwBzy7R/xoEJI+yfpwcBvqMS70iMkll0jYk0B+AiqJDCtJA0eZfYc9tTqVFcs3+io/
i6Ju9M2vpJ9Dsj0pbOPlLqtqKLOx0TmyahXUE29iZu5dI+YHC+/FilBBLXlmZeABhF0M5E0Pw25G
BXtjN5aJTeU7KgEFwfiHdf/M4ct0kxCtIy6CpA9w1FAb7UnbY1pd/9XpbGYz88vxK1ph56x1Nvxd
zfpy1Ef0XKLKutnJb4I65KJ1mTMUQznkSsERNz79ulZQDoR0WlTIMiknPzv2/diKv1NPawdpJv5A
Smp6xXLPhA20wcDcaN+BZyS8zkYCQG1Asv0i/SVptvL27kBG9Kuq0h4zhSIPwiPxMB+Af4jRAloz
v3RxcQAnVHNrkMpiDukM5ZkA6dITQy2xvpxcVGnXRG+cuk9kKqesHhbP8Ny6xiOlcVbi0eBOCj0l
UL9VlFGf/Eue9st4ZU2T9S/yiCSssLJeSoZgzqMn5HkKF/U1Ct9jo/09917N8roUpXfm+KhJtLFo
JC/PTJgjkvQ0aEh5puQRBiRObgMeqBYsCYKWDzjXRkhPNC/DFnvUclMiB9D8cDPBMSMZW4KNlzY9
nASFIcihFL7szKSXeHFgfE4+JV4Nf7A7kHfT6/iZ6HkJVewUu9Y6vshZmP1nTXN2i3mVa4R8ygcb
yl0Af2holQfw7MMwhJP+qX/L4rZNr9s/WhDQIvoU+nFI6ThQomKrz9TfTxf8qqWpj8lQ3EVtzuPi
/iMjidfctBdgKtQZDKJl7DaBEcD/3vVaMrkDojQ6Jf3OBfZq8PB471f0g2ary11oKrwLpvKuuzac
3JVsnzLOaAnbFOfbzvuFQ681/PJs1nTfrqxC+Bjxiu5nsjnH+tRY/cWMVYbSw1rYA0H6qoQOgjHo
7DJci/+gywo8dIdO0xyeBjgcCLPZlC04aavGiNVt2trCTuqgvRRi39afV0gtyS9POTdDwRSmwN+E
8BBNurEpOCl6m/nEpSSXOtOcmDHs/oUd8Sl5PA6UhT2yLdXxYH3LjJUypzoWW6wQp11uXpfv/coE
Fh3yNSHx0phgLov3HvRl0WIUJRPrf5yhCbEpZHBvSC2y/DIMaoEcGguwURLbAA+gQov93o4YHb4n
V99d8NioPSMxHxB6IgoJAf7ua4D/V91bbqxFUIFYaciDeeBPlcxXdpu1arhAh3oSXpItMjF0F8a9
29237Z8RR0lr58l6T0Y96AqSEIbczk4l3y4wWIT38mxb8E++eaLlrIu/nXfgIVWIYxnoQk795uU3
f0VZFXKIEndPXBdsx3tb5r3ST0js+ElI1d6Sw/lY3AsHOYHsFll83wON8tvquzigUJe2Kksjsfxc
7kqy5zCXJ3XWcTrUW7U6NY4IN96PuZnAqIeu4HUVC0fnJd1/gwGwg0YRK1PV3SWs69zVhYYUSp8Y
ofvQnXJdwWSTlNVSTkp9lT7KBR1sCv+mYDyaXO0KRRvUN5FlH25Yw090MDNxBgS6tysfREdykzqD
w1/7c/cXmEjANYtBR3Xn8VEtY9EYlG7qLQj+23sM3Z3EAfjHRkKaIDhSqXuC58iZnb13NpsdKT5t
OwNdKA8q89jGB6/qks674VTd3QiCr/qL4+UGMjbmgnVKsJSG48xgsm7MS6sXD6nNE0kc8/FmIrZ2
FaZsFLbAqfPHovX7q2lk+Tn37qQAY5NPG3LUhIIQ8B+3INDKl9Km3TMyAe/1FBm+nkLupU6BrXfi
2vPdoIWziFk+TvATiXbGytHRhJyrsVspAROKJ6BWv0tl4wOxlelaIsJVVYdckGHY7FXNxVWTz4gW
ZQ4Dp69vGKGmpv4+K7GfDjBJX66C4EAHDEDBnOdea60oyP7gMaa/tfWNVaL1+9NTn7R+EWo/KD0M
MI5NccDrthSNyaq+GyhmLCceL9mpUwWqqdQPLDEw25RDD0QE1IrnjNNNUSutAeY1AG7tXtMPpYW+
FNZz5N0pVKEHY75yFH/XjSfe11eqZsuu7PcoTagTBNikKBvu4aW/RBmnUpL2PFaWfHJ6VZGIxkK2
VDW/hZIcBILg8jfchC+RffQ8DsY1ftQXhvhzRl+pFkVMKKZnepszIWwvspwWquZyITDmT13axHUY
n0TqL4MG/ruuvXqOd3WSHWbxPellX2dDQ6sQvcYVyCJHBiDHEoXlgNNfcAwXXw4PpdD0FplmeXs5
nVojYFCr5UaSx72yfn2O7PXdvpmjP6IXe6NXdyek25+AW/uTuxYg+mAfyan7O50HO95s6vqaouje
fpiG3ERrqUwurXo862t0h3G4pmIUTXENuPQNVo4qtg4bUoRZBlBblJ4Xs/3OY7ZYa6Fm5zSymBWK
zFQGhKhxHVyS0wZdRv3kn6yLwzIqaui5PwltBZ8aRwIphSoanlHK43RpeLHfzePbO7is/0Ia0P4E
P4aM/Cg0AYvqWdHjhJj7wq49meAQkvQIIhZD1wMQ2dsVzjM/2wHo3PnzBx6Iw2wkHfiMAJWqGwx/
4rJkrme/5DjrEOXYrcp5mqINCfm7FJRZlbbh2RqNKzEvZRNIBYQhAgsouUPDDdN53RjuTRVlAQlL
xbcTond3rCTTXSP6d88HoUgskPjF8b5kYaKktWacZ+O2pw3l417BOTgsNmqxPy8HWg6hw8nt+PcH
+i9/nq9q6mkucPiEjHPLL4r5NCPvOJ3ycKCyJQ+C0LBP2ZAsJBGHSc3aJxRz6Q5VZ/zKcu7AOaPb
jH8lWKdttiNyliU1nsEriKDQgA3u2b68PK+Og7MSUDi4+rcvvAYzJNuVkvikF3/l915LVvf6KCJ7
Xy8iqCZljzZHha2F1bfdjkwMjf3gI1MDikpu44iPd3/NpQi/FdbzGp/WVSn8HBvLKcKAmdKPUVo3
RvrUjg6efqavGjm4yCybOIpVpCXIik5liKQToYBtj/4Lh3JfkZIGxatSogAuyKgFw6/S1f9kvJhT
PUGxeQfr9Mgc4fE+jfVYJvsHsbnZSzNwVdET1Q18Lvi+OP2XR67G4cwpLg/zMSSKPjtS41sq9giR
9vh05SLdms0vw/cHWFlCnq3jynEvHYN3JHVVgd+flpAnO/A5KBGtDezLvUop1B9g1oq9zzvIMIiP
gkFamB8h0hdU9vadN4RZMphajLFBMYA3s15dTevRMDAc8hahxmqAMb/Skdj52lLiwxOfqWt26CBo
Pv5Bb/DLj0jMyh/RvnAeP1/D5qXy+efW2idn2V5qWLqf4Gzi3Kf8uFs/fVa/2ROTFOp4HoqrmhHx
V2dTUYEjKEIYa0AmBqOG9xT0uUrSvMEJ6lo1y0rbZD6fQO7qwFdXqfg1Rojd+7v8v77lb76mZPi2
m+F5YmnKjur3H2DW99Asat+G4MKtNMxhLodUbbkMW8xUVpa2OvG4w9q691Iv230ceo0ih3yiaC4p
tRbs5CWI75yfOolCfm263zYLRDCPvdcYnAe0NMOueRaXEIDGfJCEN58/ehL8S9+jvMvU3HuVi25f
wwwDOAUCMy3kQuHR3edsL2FXfIuB0BeNVBA+7L7r9EUEidxM1CEBpuwK4pktYHtbCTaiuFK4tEct
C+vJcFhWVdJPAr3ArtQd0OF5r/YfYuwVY4dtGmBxbR/po+t5eu/w6NOHNvh/u5kOOTGKpDseMt9A
HN41wYn5PqqWt5p5zWM0rl4StO22RwNs5nGeUsk7N8nTn69dlovQNgegyySA0T9f9zxqteXrAhrW
ohrELAM7SFbIoI8muIIHxuCVYgFWBJp6LSYx07lpbtS5YRYrHXlFLLzCCZoahI3YcNi/OJrguod5
mQdWqY5WVpoaAIOjbX6zxqNfPwv7l4jXOlPvampzCUN2V9GR5G61oHtbla/s36B96Erir7E3s8dT
qOCcqZoS1s8duK+7L3PPNDF0jcE7LdhgPry5/F+O4AW64nFT6p3XiyPcMBDxqkftOSRnfqFiFj9B
9+3ly4i/xgUP8gdVY8tSjjZk08wEPPPemU7aZ8sGHjsxbuIZiBTbuB0aUry1vnWGQvIuDj27llh4
gwUN3GS06Q0MZ6K+OgwLNQyL70bZ+Vv8H/tQ+iop/ZcFsCq01UX89gwhz8w3T9UvxIkYk8pdFnza
CAYHB4/dPenJhNbXhYumI4qL3cucc3SVqmhFNwF29mgND23U67kxQ75K4AT5bW8QDwEx0ibQZlJO
gjLl1Cb/fq4vk+XlrX819J5agR4Ns4xKVUUYNejmF0wLS2imPdHyb4BsMRgyLCgA/lX7yTi2E4UP
rRl9poXwv9A6uAdXaw5AM+ce7VBtpNjFRk1cuPEiyh0g68G3epcpGQfIVHtJd/F+yrZZHtEntX43
/8YRRCFL6dFPCa58NE4jhfuOOj1NsxUHgIAVKE9yr86+0X6KDoex+oeOgIG7P0C5TmeGc12PCt3Q
xTPs72j1oHlVUswK2Xrp5IrnHFIEFlTP6+6NuwA5Cxjjv9ukQBjRpL6qGJl+YcdHFeJbBvOa+0Fl
jvNVHg/pfZQDGrQrmWbCvCq8rD1sDyJQEgcPQwQPBqS8LKdrpdoMjtqslnoxxWkp7E0+0mmuwD2S
MZ2cIfpTTllo2dfA4TtTkZK8KL1rWOpNPmrzrHtcS2YchKsjlr1JIIRHeykLvj3FQqOz2PGivjRd
q/enQ2XSiw3hwPFHXJO/VzGoK2jsiRx30cXpl5WqtWQ7H8k560awIi4+Fj+LlcHzt+VC8BFVKET/
PRcmgl/CdHcJ07I6BFLIJsAnt9PyfmzRDIjRQU8Uxlquryvaqwdltb14pp6omvghESowftmxsOiH
fQ6aS6NNDvo1ebtorymbHqoFfV9uCfRiJkwKSHADxu+Y9EhGo2TyjH1PCU3W/zw5wrv79lYiAV5k
lpWSNJjW3IiV8mlI7QFC0kTyucqnJEMvzU9RuZ9XQ+F5lOxLw5XVVlS4zz0oS/9dnOMZ+Ve458NU
b2MUhGlrnvlWKLScqJl8FoWoZa0r1bPmgO5KlOysGrhNPcnUEHId6tQt09HP8J5A+idx1tljnDQI
c5Db7l6q5O4H/bvHnoFi0JthDMD4r1HwQ+DZBdMrldHu1FJV35bD9r2PUXcNE1zqhYdZF/Csf2Rb
PCQiin64Hd1FYb7QrHY3R28XKQPzBURg44ec5wvyAPk17/0jmtNXpzihIYb1wuxVlr5rcfonF86T
oDuOKnF0cVZxpu3W6FwyM1QXAw1hvxbIXbv7Uul6bNV++joyL/UoWV8JvY/Sskse7PALeFRKbdzm
40SSL3zrnmtSa4MP1d28vo2du7nWnUeP9aemhxXv3NXvb+MwYqn1HszwTbz8nm2uGTqk7fV2feYy
HIxlnXriwx97f+uOOrXn0hocsjzngKa7fe5aljbuzS+Ve3TBJGHr1IPVgWJdpkw7E+kwvzd3Qu6w
4sQYr4yKj2RuiyzsPJzV/jSxzCgiCsOoggsIF0jeZoSMBrhl+6NFLAyeJz5kiX/Ag9sg8fgPnvnw
YOchokey6LKIZ+sH+Gp4gqJghAaPxe/TvnIYJAQAYrIhDGrXw76TkdJ832gONPswJdjx1LJa/Hd7
xBTOnAFA+s2QSeYl2fj+LqC2fyn/ggLf00UdA6KlwhABtweg27JiyG62GfdniCTn1vS/x19sIFof
+/glEALyfvMmA3qSBzVc8G2WWDF1kFYn1QDBLNnSevuDUnIpGN16jZ4Y5dd3Xcvz4KUl/cmFuAYt
I4Y/9bk1HUbowc8TjNeEbfE4il5We4ErRA+XHIR7uGyGSom0vsjd/A1ye2ltU1+zPPInRg4hvN8w
gvYDs+zMUgqr5k3o+i4F1NN7HY68fbUahXCKL0BwYRVdz8lBHf0o0qcvVg9/p2Vn13yAd7vDVuN2
8GJytfsaXgrpWpS85zxmhzE6c5jX2WIPuuJMLytnlrMowDlraKfpOhAkj0AYGEPmh3dZ7vGLTsp7
Fm2QOxCNH67UIc2IHtZ7wMM84x9S4Q7h2jzOO00YKrsIGkVTUoDJJQB5JhOOa/7uVZUKD5pspE5E
b7odTbPjcQdEbnlyAuA9cLARfmx2acYkkVUDWQdghDgxXPsOC9Ef1mm7jfFQ06kgeDWpKFPJW0dA
iyBvEs5WRiUttuyhiv4hAwZVzGkw8j0j0DYdroRPITMtcjJrieW/GI1WPO5xC+Yy5dZBc3a1Z6vI
iaplJxGrmo8RVzF837oAKSPBYvpsbropYVyLJ/e/WhhXzm+qDIeCSD1qxLB4k09R/CURqbnOCemK
rj/INUJ5s4HuA6yirCbmfRvZieKVnWhQ39F1ZGOcNb74PZIjwVyW7Mj9l5aZmEy756Ylci0PsV7h
G0x3IT1bebA+MN/4IGS7Io9V6lBjUiyvksUIjuO4VYQYVrFWA1sLu31aqYpEXLf5A0tMSfaEgTqQ
GsbhbS0ps5TIdCUsdc4fuo7t0qNZROj1F2ksPe9a0elpz0GKuxNWkOiEf7xSIHE7J4mTMmS3IbJH
jxsjSJU7PXyCtsjIYNhdb8jf4SwfIXLzGr9DNg05lQe8VClmONuUSs956H3yZYidUj0Afk7hVy6c
gzzIWn9SuK477I73Ti+GnmQ/Pdx9QJML4+tHxuM/O8mOjxi4LeFxj8IiT/++pGJMo0aIy9oggGdO
G6papLr1YfmrwLyonNtim4OpGa5R7lrEDXy9pADWCLXCHqg7UUCd0pQAlfcK3xLAFHqL6m5N2/EI
QSJCHkzIVlL07huasN3X+t4HhKwCEN7LYAg4+34aG2zwPQYfMHnxBkhjeClkI+CM1BdCVz0rAX0e
4KHTIAODXX3CPv11ykVfCOOGl9qRDfzUuLCdKIES/j1mIlef6Dd25XJrvgfPYWrMDk821tGBMNaQ
BK8CNX3Ej1LkblDTt7UuIM8z/uqvCH44hum2f6CLUJRI3aEJKtn6TRqmDHwt3HPZzTqZKioPB1hr
/apguGdLDAXgS/RXtrl8MS21Kz3QwEn1f3YHxi6Ult8smhkDA/O3RAECMbHMsHJEeOeLx9avlXKZ
2UmDhNUGhhazGWme+b6xByc9c2TsIHmeWy606DWKr3/hdgqPtZQ60NCfSbWDs7gjjR5UoczOB47f
qdHrhEYOFXNZnBxLjDbZ1Ig3cXA6WCW4o3EPAOGmf6umCcZSTjdQjAf/dRm8pchYDPlI+qUod/fr
h5SG/tTva3+d8bABZnIJL5if+3a4FTXTv/tteSlMp5i3YfUJME4NMwCL/XFKrKYfMCiGGgPATlT9
Kir3eBiyMlRuO+6cQVN3K04e1qZbmS4HgsI1DcjhGHVdX1rhDV0eZ4jHj1v4YqQCBqbcft8ypSKc
SucYr9DDsChLHs/RsLW1phct4yXyj5Xa/crSfBDpXk5esiMQClDHoOff6MbI1rGBLqxUk0DUSJbv
ZNUO35OGe8ABuZeGbDyDD6E3A4p0dDVRMMeOci3Prykc82IcSIW29QrHghkjrkcrqUgSx1ZgUUf8
/YcRwwXmEQy6G8WBjhEeNOoKbFxr9KsLhITFKlRlx6WV5Cr8eGj+2tZsnbLmyf5b5aWkiBJDhJCV
EXhwnEW/9G+4i/jB2QDKDSoiWPnWr8UV0s9jQc0nnByxiZnDj7S4eLHyTQUHYQqMtbqt3WVtV3GX
C3tfilaynu5i7k+1FX9SOg3zYAIWp5OUXNBLJbGpBMiaFdZDArbOQ//gXBFqnaPQ5jciCvuuDOK5
D4NIyekXm97Z5OHLdXsP/ESMToeI1rXWNoHPhr+0cYtXlo4AvVWbEzTpkzxXHhg9yuZVWA1L8/Wj
sEBuRPrvQh7ZqVUDzL19dnEVWqBc31rREY375WrGZFoJ9lUysOCj8/2xFHwzW1kOqPT8l9D25Pp2
nP7ekrqqbCfvl3ftwJXF0owUv5DBmdxHEvwKLUhvmQJl8lnfGZUTM9XBxfsl7oWcrHbDsF0TJX6L
vbgYAi616ocwfWaKXOiFBFTavXX9KFcHQpjFIQpGd0DXPkD6I6ew0XNvS9gVqicnIAkdrmZAQ3Sg
xBTjbUlJupTlpDRk7viTM35EbXM+EhBin80WMly7JE/kqwGDberiMko/N3QMPvSjbdf86s7M3yuj
AJdx9mi1AaMSM8jn0eBEDorigBtd1nCJhFqz4X30vNZz5B6egfEMQZPl2Qs9fF7u+yVC7cWsV+/+
V94h0oNC/SOxMYVd1Lz78BGFJokIHdy9jtftYZlAyJ3pa6dU3KPHgtRhPGsfirtBlKRLYalGuucN
hCR3q+ZKpFxGC88OSbRPSPpXDoXUuieGdudKa5KOUEPz+8aTHwTCfJiJENv9SrT79kpXKYtduBrI
ZSTqaBl1Z9OL/nuJz9cmombX3G/Gkih/zHTjGmN4IIcs7uyx0lGAc+ZFBIJjnRuG7rU1nUkw7yPo
QGqQqh0BxzBYftnQRlyYkC30r8XdddInhX6pNEHcF9Kw3WKTkkhk5CndMWhdetL+AyTzKJHU0RUn
GQNvpnwrHFWQ84NGVkJyF1NUdYqMdy+bXONFKXQ0sKhMs3pdHsYlI3bHQnSxODgNKC75h0U8P/Nb
H1PxtDLcVzg3Bwa9o5BJTPp7sR+c/j/l71Y9Ku6wkN7OZBfqHWBPZitEU/W3t8kRxIy3Rbzb0aI3
PaXTzmL73iYaqVL17cLvpZwiRZH0K/bcakCa1NPz7spsBUAuUfkWnE9IdnnDqfvz60tmruCyjRrE
IIGwEZJ/Rn0o61fh1yV9mdPZZk4t3DSD1GQyjvUCOVsxYnI26oB85Ssbc5/HLRxNicQhywfwH/f0
zNAlYC0yPfc8XgeHg4SJPx9T6/z6QwrW+NgIp1MCV0uwqJvtY99WEbPbxmT2Bevcj6IGV75i0rrs
sDhtcmW6c83w0MgZUJPSMdog0CDu1PvYDQATA+xYZLiUnQxu186BR27WbCFjyzbACH+eiKPzevCP
5Jb3y5KJQuyGnO81D+q6ZqWWDayesUG7Ww5JttNrLnGoiSa4wfR/gBrzPhUd6iY3Ixe10JucQQEB
zCu65AX9u1q17LqKufW0J6vc6BfzwiGNmPYiKfND3dk16NRYTVT9Rxj0Zu5v/KgQ7O5Kcho81Odx
bHTANVS+UGNyxWpD80sYSIaCHemuIccEHAcqBrOpQnME5cdZWWHC0+QW9gkrFBMpLtwF+bY5Gr4W
IiyEDy4UXd+2s4HWDZtVIeym94BntvRABssM33XWpp4U7TlHLDz8gsEX+dELtOC4LgWyHiY6FFYE
v1fbMnsQOfkuPb9OuK+WXG+woGb8/jDmXinn2vAq6AzKwtg9vht8ugJVfye8WQeKPsuNeH88xKlm
aVRJGD9gW2W4fsJ3Gyd7bBMtgTfEqvXDWWUEBzyjSMDDSV+mhNlE6M4HIQmWA6sbL/X52ptwPN0s
+iF5bGZI4Xxv+BqOStWNYS+7AYFeboTXZQ/GU8odxdoyITfDws2G+ZToxqbKjDpOwQFCiuBVO++u
yvc0ee0B9aL6A6v4oJXdy3YpVwTD6eih37YnxT3dH9ImOX1KW3p0QIXjY6t4+MqP0PpxvQKVUojt
bwftj0nGoXW9QmNsdeC/OOgNkD45+HHNuImfNCYAvEihpeJ30LkNLnNEncrhpZh681m4ds7UEUiv
EA9SphFRJnq+SBDwhyXtZD/YJhmE4rq/zNwDjZPNI++UbWUHJZxb77x9o5WAq+N89KxEF4eTCHsE
OJCd0Di4BkCuptyEHwZEA8vuVeRc7OMMojdqXvEUJbh0SYvr/jGrZC8swACdFdXbA+fgtsFTorgJ
DPgfXExu5iAr1No8XNeYGGUiVP3TlbhhD9QN5y/b6y0tin+061keAJ9SF2Gg6pEjJhzdlQ4SYkn4
BgsFAvnm7nBqB069NAkEwtJzpy4h0dDugmebtELImDcGETfwU/uou8Vjj18Wyutwwb3oJ2bTUtpj
xbHdYy3ODfuf/BpLN7OrOcKGQKvgmkm8fetO5+Av42ISIZcrIRDkbZ4h2lqI6V3MPK6VKvmCpJlK
eZaXV+UceQ5mxbcqigsjoc+kGDMitgkSVwY7x2Lvru0V90oSPkocVmfg6hwh9ruUwtsSb18xyc+I
dHPHAW7ptb82SgYn+8TXATFZn5aWqciCEXwd3qVJ23HcCK5CoKn8kS4kFYqqs/uZ5sYJHsITKzgw
87unXH1jeWiyjJ75SUUzIYJsyJML2mtaGycNNf27DGwT4x3vIuum7v9VrFeY9vqxxgYoX/3LJGv5
iJ4e2xiOlGJN1/ELKdh0n+6f1HGgu8RUuW8Ff101vLuJ6kWsbsh6d/zeoeK67GYtazrluUw2lbyy
sxz2h4UdT7iPHmgpYKuW8SnZkjYMuofgDNGKQf32LCJk4sfdFPHJmaalylHdgqec3svjidvTknk6
+++yg42537rJm+iWds0JBaKiwDM9G/TLiaX63qulSS5pQT7LbJpUyjW2NHY4Fwl2YxlhXohAqGdh
4QqfbYciedxrUleLjMHOSLB0VEVntfFXmU5ASkKTl0iEpZc75oZxSg3uabcb46muwanPrK+l8d+f
WhMFIzpZbosXwSbBEHVi0cBS/Khd/8crwiHVaei+J+Iatw4hJC6NH00sT26ngy0weLY+U76l8uSI
P1ixU1kOjY1cZOq1UjJ1Sa2dl/aNCzRVEZMwvc2KVm5vq+BSBKfj8iANazq1Ol0fSwn1Q8LeHMqb
UFYN9EID4BGn+q6LkA7MsDHBA8WBwwaGfR0iJf5ih+yv5TvvJUdU87gSP+fpx2jhU+6LoLqB+652
vr8cGi7aftFPHjcuOLap2e+jMgup7p77t/rYgVoD3j1pYTHC7PhvSvl9ktPz+kmxwe4Zd1veLVa5
0Jny4L1FOHGMsv5u+E8bse+9vxw96bYaADvMbJmkoIjeZKXRhoeSRoBCDkSTtFIb4Lc0yUVa06JQ
1DPIR2YEEJfviYnkoItgvvOXz82qpM3RLhFQRmE10ADWuT5nG0avqkvOZH9ctTTf7m0b4hwkwbj1
UXGfnBaXmLWv7dO+jWcyaiemUfhZ9VYA+mdXNc/f0iL/sZMLiQrJ7yofFHPUeiAZ3TtM6sm0t7zc
owrgVFVXc6KjnPOj0HgxmS0zNU+hOXmgvs99fFBwHP6FLQDrWSqDI3IY9jryA64WSwpeDLe/SCJY
GXY8KZWWKGHZPKSpZnayQ+V4Zsn3Chn/K+Fdd8itoCnyae6LSatiPBxJl1nfY4jOU5Py1Y71DcFd
RPYu8orQQhV0u6/HWiPxZd05gxUYLf31xvq5UEctEwSVEdkTfH5YL6KrxhCtdQoM0ZSCpoq/a6Fh
rgnwVoIaDMJQYEL32xt1MjQG4183OV5x1s9s628yDNPULHI1OFt9UPMnROVgruI9P7fxh0LtN0Lg
pzNj/KtsVd1M0kbF22UGgdjjwiuKCldvTXaN1ioDzWI4LCoj0c1kS9Utl+tCTClrZUxeDt0iDjSJ
MrRQ1pGrJP5e4cVjdaaAvD7FDhWsJpMPk0iyZVZpjqqG10iSKESsWocvrkYR3v9sNJ3ifJtIyvT/
GxBXjY5YfKwzHAfDXhiTbzrOWmK20G/1NzuhF0w8iN4HpHAHPBJ+pG2fYVJtPRqn5wNUSw6rcd6b
20JVcth2WrUeDRg3OVZ6eQTEPzyPSw1ZijX9tfB64E4IGTQxGMGk2fSSll4249RD2laD3GQlKl3Z
+nrq7J26Qk3uahZkWxD8lQsN1kKBR4Ul9NXUf+jdh48nx9G417lfYsfNyMbwnxwA4UquPelErAp2
0niZfP3DTzTdIE/zqMjcMcV4eZCFaiLazEhkiOAZjXVCAvUEftj562mRL6Z98cAxBC8zmFRNrrWR
D86ln0NJWt5ofAneSsWQ8oRvhPArpvW/MEXwmnQ/JUf2+G1rRxpcqoielkwfhQHh3KLfy+iUDyKK
4/C+/0GsndeeaNyZFroFa2fhSXhTb2ENjynyYQ2a47kxixd5d7e8jcBYnnEXag9ZM4FzVbn3nHmF
v/u9li9KF0adAj90nsaxYChouaEU8WvXU1QL9x+7sB5YKKWjhJuoppUC7Lpmr5PStfXULAl/pl5U
GzhKfB6qcDonSYuilMriyd+//en/26GLmzgFHglHW0Z3PkrfcNbaH3zMH5ZEAG0/qbzJE4biNNtz
Ll/qqk9vfHyIXiXwZ11dJgumVCfphMKkU152MiiTlhSSCzUoWOQF7iyP7sbXAqhI4si5u0DF6JI2
yznwpfgTfzqXAVo503Jo5bIAI/YkiaWSIy/zDyK5iU3jen7uZ6ymBOdG/TDoRVIVkPgwFaPih/3p
ClIpDVT+m0Sn+H7z+svZGOXkowQjXAfeGtFdAL/zAyU2O/Q0eks4LDd3LmE+P6vidvhSiB9I2rUI
+9WI1+yCrduc8n1jImXKqBCRKUW/5YkkBa8zW3m2Zc7r/jkcEmg4A3R5txEWazzb3rDFVNcbdGol
+wjf4laFElbGnthbM9Rvg+QUZWZzIf8vyWoS8tWe/c8Sn0tY9l27upUjKsN9F7okxEd2zv+BS07x
X8tGUN7WmK83vlNCZwKAOJjlGcxBcxylYgcUtTvfQxzik5BlrocvyStdSlJxRPxXmgT+LXLP5Avq
cydRKimaEIiepOmNpJ5zdSc3q6eEhmHa5j1HmM7skol7Oblg/Hb14vyFeWc255hkWLLlGS6AY56O
fA36QGVRSyve+bZa9yW7XH+bJX4sMn0vkYPnDlKYYo9ZoLBUfX9tZOetj1+nkJWrLdIZ/PwsmUP4
sXB25aBOuIfnevJocTYP44jjkAtbZIcrqwP1/c12H5o5Blauu8bqqgLRllUORiqF80ttXFNY7P0v
uE1ek+caj+jUust2vABUKHkxSZKVL204ZWBlbPsIMAQcHsjPRCH05O6R+GBCjJSnIMQEnmkH190j
HbFhOgJvucBga04VeJaLhZJFe9yZS1xrmu22uk1jYA010kguf1Wfr248mUCqHiXYJt3Bar+aFWJk
mERA+CL5LEs10h5Tl7Ajo4yV34n5kqrb+RlMHCyNn0Sd/USRZooymxy6mE+RO182l4g0aGKq45H2
UQcBl6WEEgnYc5r3tk00Ii9osIjh14b5uMRAWDqitZhlzMUBlNn+VB46BnSf/N9EjQeJ1qK4pvZW
bzzIVhfjcSBREHrY2zcXiNvvOhVa/bwUFEnMKOv3Cf67QQ6p8e+Zagl9RfR5P+JHeQToZdcf4xUO
hQh6Mxm8u58OtafK9Rw1BL1sCN3lYem6gLM2LJCEtMbJ2OQqSbTET0wT9EHDQWLK+XpPVCJPt3MQ
5jD5PXgyg+DlpUsrCGyiFeD777wfRnkgMgM5OaoHca//cYbDND/wJLpCveNrRjQow7+0c9VY2NYu
HKXjrEjYs43ODwGujLEaHyWc+Tonmi4uO2AZtMTSlNlEw5VRlgsd8YS3r57s2N9kG6xd8YFeMP++
qs9SKqi2XdDA74xr711OILxyaXTWgTAmeFim5wXvzG1I8kaFo0zpFNFEMpe7fJ7kY+tJhiqGQFCl
IayRBmmTxpW3eW9hkE7Ez15JQRiV+CAVhfxKw/2QbpMp1IUwxquksb9SNCVIVgy6ciqh48AIM7ZG
iLQ3eIpLbBEqPxWElo3YlClnORCS87zgfgYp5fXrGrxNpnkfi82DR/PEcAxsgcVbuZi786g1zObo
2n6Eqe9HYDNaLNLKV7G0Zf22HOkL6VWIYJMvdZAZucX9SYSjbZ4KAgFhmNltjVTMfyBMZaZbl8i5
S4Pg0md46XYidfLr1JSm6X7CDWvsJYcxFPgQUm3Uxlp1L8vheuBplOFFC7FmNF3uuSBh3Z/EN/rt
e38Sb2HROMqCrAPtGeZm1RfWXfQjFT6WI43SrysCtJJSJMoSyGX2zFNvxYXT5mltlhTCKrbepTsC
Fond+pEfidTkgzPgGVzaLpchTApG1RjM/R/HJCWlEEaHu0RfUoegbYatIkCHSsgyq1OUzw3Senp3
hX583Nfmi7e3PHPp1j8kyM3maMxFzuv2okUHexGINYaHoni795fHZHIwxq/FtMlsTJPy8C6ZdgsW
K/AfjbAF1P5wA0JjeNORwGzEHSxYWJCQKiRWoINAGARdwh1uHCcS/Wxpd/xrWREkAJqVcduEddKj
cZEJ7ZE5UhL5fkGY3+SARuSAmdze0bRCHDw3ilTWomE8RT8Gh99fY97gqu0z79ZOsrpicawkgoZv
yp1Pdz00YU8Z2xMRnxDL63S82lPwYPN5DJb/7yD8+OgrQ7CLDgfaeWG40Poi2b+X/emRwOBRaq1O
c5wXrn19Xj+F0UynM6q6lr+Sm/wlfERGdMsCwqTYM18v8DjVFGqzI+nGIYxX4k3nruufGX/i9OPe
l0QnkKpUYS6nsSVPQtN+QsG7PpG2XayAPk9Apler8rd9hsBd+ILjy6jkcwJoQbVuoEXT2sOO+FJ3
2sntfVn+IPwE7sDfgotJDn1GBYmb+aAcMjs15F69An/UqFgIPobsP8xgac6KOFv8Pud8powAVD86
hcKZ/9mOYhZvuihEczbH9xW/dqxtmGmCLPncfc9JgfPOx6ypF6dPLtiqC237s6ZLDsI/D+GIldTW
OhbTK+br2QYBgFrpXN9UPr0leuoJDPI/VKyU3YcdQsYPmJKoa3Fy3FlZ797lIWPWNnPLAFcf0mCF
lxooh/V4dl3FymWeGriNsiKBsww4yHodeSxkFXUJDS9sDvp3Sf5cwFvmHwcrHGa/vL/87G4QX0Ny
MujMHfFLA0tXu6JeJ4T2scTVtcDBWrzUeTLAAFUSpPCSIubE645D0Z7d6T8IHelr+YuqBzQjYkUP
wDTHI7Bv6uNmh8+ox/b9eVYQEmY2F8H+HEt2hNr2pSi5yJ3MmJ7c4QTmgistbQUALgwG34oJ7Cz8
8/XUJXsHIJRbv5rmBLrqQGoW54ITKBEYhJ7HVrI/bEa2zDBLtxH1WQGQG1dB2Jc5RyI7ji6BfZZS
zja25kHeHe19gFfidb/HymdzBJ5vZbQRDYVOD+7dRgB+DosEbS0iG5aH2tdUF2GV1qHjsmyRax+l
6FUOCbScNkJq0UX+EDolqo61kOm5NUk+OkHiTqABC87T7ghDt5J1IskGdzG4j2vgdd2wnyx/vnXK
9G4gMCZZQgMgIG0fvn4FkCwNbYUqyk8Cd4Xteuy4WryQ3AamYS7fO8/kmOeJGicH9zfPSSv5W3HC
biQReXcK6Zpql2L9a44UUlkpXy5mvx+aJ5GIT444DRPnsBCuBAY6ndp4yBt+MwXm6oeWHgrvusZh
pbnGqJNbyjUDfXLsct1DnfkvROb/Tgvsas+zGXtq6icUy1XjuKd30bfithDML3lnYp3QHO8gxwVY
wArWUjdCyb3Rh2OQ1lW/XqOJwGe9bu/ULcWu8fLKw8j0NGPnreox/5GRtCErqW5XPStQIngSJVuT
OVrLgw8s1HeEYm7BSgrm48bFogV12eO5PuI/ol6+oStyjwbDbtUBuwjJHU1YhzsRTxVbTMNAtOP5
iASFTnyMhFQhhpMn++l14PqO0asBsbkbIzNEoEvTcGU42NnIn2SY801k3eASd03k/vvfFr1F64VR
PSAkLdo5PUiN5/OlGxsQYt3JWpuY66Vcl7NLsc/bmdp1xZGMPjiU8XRYCadXL0EMJWvvmpfeK9oJ
EarteN5wMBXXeu1NPNeiAaDz+pMxZFGvrJAaYRsvhBMFRnqhtOSpd1NlydFoM5zih2IsAuzy+WkP
1KClx/+FG6noW65QStfIYK6xSRp70OoDz1Khs4jlqnbwoRQmRLzr4wUeIsQgEwdAQAhcA4RGLLpC
Uo1Hn53hLHOez3zjzSfwS9NI5I05kJtFyvNRW6QAzDsK3/loNT1CcyVdJ9Ym9KZbHxtA3m9dicSE
MqF9EuV3B7QtPJJc6Z5O6RQf77+c6sF2eEOKu2iKYP7FTcNJeXqvYW0GuOP7bKZXZe+2bunpf0vh
DYQvSI1Gj4zhWZt0WJN7ImPnG5Fmo2pzFBPDqHbnpETqF+uvTB1w5jNB7HYKXYrc/0s3OrwTWo5f
7OpSI0v2+Gta1/aWSAtv+DmLmIxEpF5EL4svOztgZyWmGda0mwBgIxU8qGHkNGPXjgwcZITyq/pX
txuR+h1UJRZP73A/vJtPy1nZ20/rRrqMu0D/r+5d62p9zryJWSa+qnZlS/nyfnMQgfLI6EXPapsj
aRbeMGs+U3kqe8IUOJ+T/GuILnoiUXeVVDs3jnjYmwWCw53l0QYjufsZXq4D8tA7EGaQtotu4MUo
ma9xvZ+JFHcsO1fmLvw2xkthBNWTiiIqsnDzUAQSzvTQJAx6CYdNAXyDjiU52a2H6DPA4sOmaoIE
YBYMa1/07oh3JUyRTxock2UU3AfVU2tcsz8j/yW0j42Pjg4TnUnW9zesBgmEeOcyRkVmcNUONL/i
Dh6L8nlh7WFn5LfOA9Zka/WFPbyTCt7NxGRlf3uCEw3WQQuK/J7ulKthHa/iWR1FamAKFGaDDMQg
YO961azjztWT/63zwFdhBiwDGdIt7+8mXpZxgA5CY8X829V4k2Gxmy4Zx4nVvUMKW/LoWdAYUpjV
zB6j7e5oJTmJJtDBzcAG5Bue9rk/Y2H73jjh+pNJOFJOK4820HjwJtvz79YzYqxr8sNZm8VPwEV3
j2Kfc8pv2vP6VVXObQwgp9Jus6wyfAjQu13e+eCa1T5M2aJqQHGMLPFyyyOI5+82FBt5k2ksw4g6
sI+P0EgQC5Ntwh5KGyEmGgaXAOQjnkuECM7bwLWTl70jtlZ06tmA7nP4dHAVMMChTYJ7C469MtHK
jxKDEolMoluBfU4Pl2mGQ9RDJcja2N4pUIktj9pA8wuATMsAlQQrBKW6yq7cGIpJMYgtegZGTymE
7yObMuqCjqNIIxL0DV5iCUqOY6nnwYkAvriUewN0QHSZ6u1GCv/HdX6Ku7BKsHje2vEieVwVpw8i
OFuPABEWdkp4ZZOIplQZJJ+RBt7kdHKpAPeblodt1Stzb/Zx0sX9MSQOxB1qUk0QW13Je8EVqKzd
NMgKgAO4bqNSUphb8bH/28yLiqV9yNcgMt3uvkzRrHhbX8PNsFvQiaZ5Js+Iu3SV4EJ7sQgsgpyM
63NjG9wFB+RLKJnvlazn4tyZ+Kch89Rw83dHB7is6QRvmftY/7PB/js7kNzorDlU0YsqHhQK/ufa
RgBxX5nGX8quZZjpwRyRN07T6JT/kuvbYYzIoPLqcrdybtRTLd2Hl4tZvQayQ6TOtMF55+aowFnQ
niNXgvyZwqzmyYm73kPSm1d48/RSsqQGTZAbbgrSTGR/rLZWxHDOIOx6kQyxw9ZQ+eTXMhRWJbdH
5Dpslqjz9ElL7978P9UAqaeM3thDkIO9bEyvTID+aQJ2bbKIfakfIGSb/gJPwnfVsEecCGDOvk3q
8zbC+B7t02E/V5EZeCk4CI9CMC+AFNXnbbKTXmhlsaeb2zc5PGjwQU98bX318LcnKR9NLVz6NYyl
1ZEA7kwUyHSphZYqattPMhvOs+htFYPdaRX5V9zkXRH6oO2nXHUmkovtq5wAYl4hbfiwzCU0FUEA
pWEekwmwuAJCGKXIzditfJTiXGGwYJbvXuupQLPP/EGlZNWCxTzXKrKWGDopriYsrdiHL5O/WGZm
UQicvUYrGJMEss+LsHPELXOY8u64CM4a5zsdzSjGAtxi67MtXaIOpxlvNzdhj92JIDPtBLKC7WWn
0LIcXRqOxp92IlfqXKQAg76y+ajOQzu+/qZN+oq6uFUCNmlwWC7G9AU5vbTg/66C+oI2HUvyVHct
fQsxh+7KbZUv3XIph3ZOJDv+9AW7T74wgP2Ss/W2T9tq01PsSSAAQc3hKEopJFflHH9K7rvxXK5d
kINuzQ8RKd2YQ5yTiIq3dwkovHin2TlHJaDL0r590fZGSNz+B683n5kvw+5/PyT2njUJXkoyaDmn
Cej1wpa6vAUbCw4kG3wtkEsDtP1APbMls+vUF7h+CJS+yhkSOlMxsfCLZnJnQ1ucypBLn4qLk66O
YJ3hAwd7rzq8/xcNaLIcAoR3KvHYcg+xLpGCzDXW4kQ2cZyV+vsvnZKXYzZsgXc/Vg7R5keQN/XQ
0e34pL/ThxcGvk2uKRTRLHgjkhl43k1PmUUtcaiuX8cv+XWRsu+FF+0Lt+dbJ3tiq5AWtHE8w6mA
+Q92vHhRjrFqZEm1DN9xZuMTgdzIDuy+rEDZDTQqt9BcCyz6CLJ25PExZLt1YbyeCOSRbEDtbdWR
VXGNUTof/71K5iu6E96WqcYPFad8VXKkl+iiFUe9gZwsnIcpuRkgk8QWsqPv8S2Qm5vVGhJGUM9N
IP+aP9eH+7Ha9jRPmN69R/Ze968sY7OIpHBLOPsC75u9ItBSx/SGNRXcS3wOZ3SUKALGXaHmvC1w
eO8Z3tVGgwO6T6Vjwg1U5SglW+0frfRtihX4w73t/PvMDY6h0hJcG0gq6SmfCu+MYBgi4WxIB5/+
FRIgw55ZZ6orB3h+JA4IanV6pYHawvnnzsjjxgslyfPr/CYv8av9bG/ZQvjiq01fXWHwJARQW/t5
OnCv/CYEa8b9EYZs11lJEPeKMxP1SOGNTH10mYFBoWclcjKm0sfmApB7ZGDQjBci1GsvL56vVgeZ
9IGYjwDO1yQU46EVsNSOZs1q2W+fwxGKLY48zg72nRdbPabkpCQKZMIl4WEas1odGIH5VfGp4jUu
hC0ebqijIogGFV/SfsQzdOsjXR/39P4HrRweIi/Mdj447ea82omvDMaL+ynzACoBRF/BqWtWgMK5
8fkVByMY2FzlS4uSe8+E9clwBchnFh/71zadyHm7l4Kwwq75842g/NHWwxpOLRPrJq5hZRSQKwRk
M59uVNjUuRUAoCyOXnci2SjbF6tq3vsPvgYNh2U4gW2elVkhdc7EICk6yApUYLM4r5KkqLaxKwVE
dc74GHaIwMyguM2Abp+64yCglHXxn36NjQhN84rxEv+UhZ6MdUpapoc9yRAiDzKA+pffvfCGl3TJ
GWunyBzl+DarR0926H6/9szXU8AXPZTRbvAIrbVQira+84/xRmpYL+1DlBKtxXoDhFahvpcAk8W2
Hc6hMhBUY/Lew2dk3xpqTi4uMJexVurPCfXHNS+MjSUAJvLuJxT88lzcShtphDDSZ44QaliYokQo
Y2GfLnKwSJdU0o7OGPLZ4ycli0Vznk0PFHUI0qDZRECw5NPf1FqRigc/9PsmNEU/zQPTVxjmVoLO
xC+OkP/n0IFVQv91FfExE6XzyPRrGxqSBW3CG4En5A7hU0+L34XALg3eN5WgYZUI3UtucttETdfA
CW6QG2G/9iwD2HHBBpfCKPDKksWj5nnYSL56ACs4o0RKUrz5mZrpBHjjEASJwXr39Nb+rVBjduim
6zNtkLtVpR2DS8EJeIkZ0N0SjMn3uyD6rXjUjbneY1SWAlDOqCCyv/zWjoreKH2zVs9T1AWhFg7u
3cgEFwfxN3vYm50Ig66Blsy5gagvthnwDvRMdsxo7ZUeCnxKuZ4AkngaT2GBUgZzzm7SvAhdSlL8
Z5R7RXQwsS/rEru+cCffeHQ38wg1LrY3k52vE1POIajZ1W2vn+bFMoqr+wKjxoGlP9cOpzhqdfkn
/6EnW2E0yEzr+teYpHsXMnWJnkJkhBQMJS9jPSRe6zIV3YVnhz3Yl3TCmsE0LZyer7GsnQ8Tm3pX
SxbWviJDyr72PABpfFP+RXYpTJmkmPKnZv6/lvRbJP5uazg4XVADD/171qCLWYgbGUJolb0hLf9L
JGxAinPOe7m3VwbpjqI55vxHy8DEENL3BVxaL37ysxENrJPdQX4SIU3yEcEzGadEaWjFyz5Zz2+w
ZAvl0xcFNwb/k3SaSwkuhopGxqmuWLvN1H3+YQb4yzSeQon7/bvxWILDB/eaG/Yxzhbr6dwKzOqp
89t3QSuudBfsKMQJ85paiGkvj8XvZkyoz2Ni0WBa66NYsK9+Yuasp+xsAW4qvF3iLZa8E2wP7wl+
8EEU5w06fOIbmADG9ANprAyKHvFBnZ6iEiIsEbVcU6L2lPzOA8l+dpBqvMO91LHvAVj1L5KrMV5u
+qU+ThWF+LwMLjvFH3cnQ6yod6oIalr01qHErBb3UvcCauWsVDVKGpHGS6BHBzMJVAgsNf/NymlB
QGCDe2Gkrn5l/A9YmTCSGY+gj1TmII2IIZhEqjYXnQ2T2bRSmlbGWqQx41TLY4sqK81Dgy64H6BE
yRooFYUBzVgNJ1ePBkq4hlquESiL5i6tFXTEldk85QwSfwE2aN1fPrZBJHM1nE/QBmV9hpsTsL9r
79DmC/XNzIaVLMVSnfTspTxrCXinqVKBgVuTqHfqmvkPo0kU09YjXDMArs28NnwEPwagRhlW+C2R
GnEyCIaTeK49eZvWHoRYHj+wHtVXTuNAZI5yyl5UnbSylxiUvcXI+raYsJ1ij4O6pMyh6/CIr6CB
uue1tdvf4dlEDJ6B2nrUkSoxjwX7dV3pxnmHyP3hRJ+yds7XXzUBNOgsALiEOiB4xtJJMLIX8mOj
I4knMiu/7vqjhGrI/qeaRKH3McTR9CWItC+W9GPWav45BZ+v9uuunHKQYsufIN6OU1IXPXa0sEJN
tmX7gBDUjiI2GNSSPpLeQWcGxGBAgjEjagimoh1ww+FAt0LIifq6m6+n0/h4S0U/VzgIh75x9m2A
Kfdm5hPHAh9zMd19g3cvjYls24yxN4r+vURjFA0fn93SkuhqMZwaeLlUVzB1dT9uaIQfogy9cSgr
h+kwE0zi+797Wh8s2kejuKk2lSpKuzYoUgVKMGhAwUm8nyfCmhZaoR4SAIoAZHBvh1EnAXH6aaxc
UyVoMTZGz9+pJsY3fqPonS33R3QWCxQwjcm1veq5vPu2GqiSNSH8aM0JmBv/8dhYYOuABNL9HGxd
j6Tk8fLgnOor6kQxrWFokoGTgMN/uoRUKtW2+U5sASfCa+PpjK66RvW4C9XS7TkYDp7P7JoMK8ou
ud95MOKLTSn0V6R86jMbV3hZYqi4FjvnLIy3i9qjsRARTeL9cHRs66OExSCqqp7LFuCnR/nAx+Do
H0X5l1046VL8mVh1+y+B2Lb0HQzPM2aZPwq5g17KLETBJ8k3ygTEyOEjKba5yzM8Mk4mbtKKM1++
cfZuRLRm2XmjadQ9A+p0zuPqO25lIFclYpVp7dbg7NBuyKObCfxIbaQP/qPtnn/88yWj2aSXLtN6
cD5bTvZyUmI13xqhIVvpL4z2JpdCVu13jb7oVUI2yA6v7mc8TsRiJc595peUnXNlHFA2LLFVkdwn
b01DHu4vyDlL5Q5ggZbZt8YSGWIgR0eGUwQshemYQ/3FJMj/O1zfVuUsHz7a/aD84AJWytp1fZlM
xFMPPfJrj1KGVCOVtVCsaTHkDNhcDxgugwFjhNUsBeC6KeA5iP4lPbUeI8DoKJ5zI/3ycyFZEzDK
Csf9RB5IV5gLWUEDbp5amoFf57lto18lk1uPoqZSk+vevMxXpcA20wpJRu7Apqgknx690RWKL/so
oiqnpHUU1J2gbWK4rB4UMnmuOru26LYjgyclY5Lzgn6KIbY3UccVGllzE236kMrAXpkVFhraUCMc
bcF3RT7NBSS+MyUsc5OyeVi7od3fvhdgsU4nwFsNC5uh9x2ck4zT9/1PSOBFDkS9mb3FW+KEmp1b
ee6dQSVhVE00Aff97H9Q3BKz6Ab50t1ls0a/MvcWtzvAAQMOpktAPL6XjSkKdSU9sre+DqXxPPZ3
6bxpKxepwU6O1RDy6+j1TYhlZuCu+EIERzvZIOreXI6IlhM2o8dL1wzZ3IcbhR5c8PXplts6qZxj
2kF7pwtsdWsc87HxhtSh+yNieRkqhDVQA2CUa4mzak7/Hhm1S0VQ/rx0fbXfjRpjNA1zukRIHl7j
VsJdiXJv95imXZy8I0bGmofjk7mdBMYokIduUEhHmE/gZgbPHL11Ifc4lvLg7AfR2XmTPfYEoflK
HzXZd359nOmEY96CXj72ILc7hUaXoDnEwCl59XasZkW+VCl/gUY1MG1guihvT7eCo5Scvs80PeTs
5TijVHYMpn9nSZiUxADVpyVb13PKoyqu98lBjCdo41zyieNj750iRLB7YIPQ85OT9zLrAB1jDQCw
8P+4U7lGvT33gcc6Qa2NvFPp7LtuH27duGDoOCRx+gGn5mG8CO7P9M18e9PIiN6jRjX19Jh+ufNo
/LCMvf9vuAAsWopVNyzfRowHiovT71jWMur+t9zN6Q2/CJqBwqi2ilwTxSVKcJ8jP9Y2fzv7ZFP4
31BzHrdE8Wvcyl7OSCJmfI5Kr8GB47gUJcF0NgP4qmdwbP0qcK+qlCXqFrO1P+ACPmPxE9QTg5y8
Wtme7wenKAsKnBMTcNnQcMKavnz8+ProWY7WQPkm/61/j9kC7M/3DRssal86NZzq+dehOtrC7PjE
3o6g64qLHijJSBAPYItnmeNGx8in56uL+MDqDof1zkSI2BsbFt4LENhD8RaVxr6krr5l7MBWqQs2
HXaYQ8xOKF6cgAbKLNUy3P+uZGvu6Red5bVl2jAjM2IbNHrv7EBfvqsJHxJkR9T1W09q1JrWRC7F
IWsmvtyTJ5+jRpsi0hZwCI89RixocE+Aa3D99gy7rPwqIZHymcJG4lT4as1Jk6tuisSG9qUnOORW
dwjfBzz/QvSaozHw1fxZ6/aAmaTk0bgCp7+64Lv3fWuAvZyVw79mc9710i/SJv5LqYk1oF7XS/jS
fe3L2RSRx5mO/0IFSuT70m3Bf2QQY1zgtho9pSrCCJq+J2jk2a3euhDjlSJnLGVHeQapDAFRuBkq
lHxrUC8kqjMwyB1OF2zQIMXgYF5bwSNECV5OjvRJQpr/XrpGqgD2eJsXZXcnrBz0S79uRA/KkAMW
oH+5n2novqfqJ13cCVxsxdA2msTge0vKiudwizCpEJiEe9tVtB6Nbb6McME8b1gIigrHhKQCL3y4
eVwf1s2RxDURizEj9bnj/7stSpqz3dUJUdNgPTuwhsflZnHEFtzR3DXN4rRDQ8Ck6PynZghogK2Y
uOb6JtSwfKVNw78EAvEsemf8XXhbB5lsVGsMneyi7/xMDl29icAfrEuOMyz8vnIyl5MKjEoD/+OI
8Y6tHEHrnnfH+ZJdda1RlqDm91zqc0i8TUCFUkgnXXTF+OIPf8YdmpeVdJCMH53P61/+lX71KZw3
FEMdANTrjWNmz/xKV0qx8G9ePRft0GlfI3qQUKljjx78Q+xKHySbd/BQWn2843VMBpiH3DiERbUJ
Uyu5UKRnuhW4ROcuoLWMqTzwwW7P9lJK1vMjd40yJhXr9C85BHdnNEBK+AcsOBRazorTIIpAhEan
sZfDhEpu3crmT/LFXWnz9ytAJC9miCO5xcrVVjA45pV81NAenMLvyfQVMELqMQM/dMrD1+Ww0qDP
UOJ225kl255h0bA1oBS8XaOYRxFdTA/heXrP/K55IGJ7m7TNNv/aL0er7J9w0DxqdYGIZT3azoIa
luMMFTMQJawVmQongU41EJhMIRE01O4SUD8U0UwfV5RuQzis/wSUa/7xjpmWpQmK2opbDawGTr3w
iJg7NdUloN9AGBPcaSoWHNpW7XdBrvdYYenqxaoM9gMdH2k/c+BOaYGwq7HnHdn8r/qUpAuhaL/n
Yyu/hh63556vGjPeIiyF7HtYforaGdFfiai3G9j/qqMXzfJnQBQgzUzQTN3Td8O9EUxfmboASOyi
zPoRNun4A8xtB2cIpYvBt+suETQ8ibA3LOwx3P9xfrGgpZUsR6vmM7M2UNRsmwH4fg1rzS5+dDYU
sbdyZaAeShXBYZnSRCfVidUBx3wo1emS/PqPubERGsetG6bdnzYLMKtgMRSFDh0+4+4KMCsX2ga0
g6TNFZGbCIIIH3KzZqkSuP1Iw+5DZX0keolpSoLkBVNXav9Br9VZalPJMVJ0ITQBnlwvwSIFnv0s
AriQVAZKNiydflBxRI7BdkCCoW/9pNL5mQ7UWS5DqRMeD+69KrJ3lUboXRaT2RqxL0iPuFpXHZ86
6x++UOlN4qxGIO5oAMxhwMVruKLNVNRlxIk6HHRQHesUBQIQaYDoB2v3vljiemFKFvR0qiuXvF+8
J03Vyn86ckZnWb/9jPgZAcPsbJfmdf/Yvau/Yfd9FXyvfywbki9nrRPJAFvRwpFIC7r+ZFUHN8br
aSo+vg8H81ESJ13ALSPKIZ+i1rRsDYne17N0NaFwtpVGyxBRQox2hbGEyyLWLNz4rNgejl/yF3j3
y6bZveA7TY3B4XH7AP1OcW5oJGaQBIQBtG/SVIk1iqmKEdT4FkXyKM4Vk0/32U9Wui/Cdlk2l0pM
nUHHuYOYWdbuSPzG9ZhwJiNTtsA4xgaJdm4RUUvjEKbOGdEyOmv5r5zlmlZ6qWh7OVIPL57K94sD
DMnUBGkUwYWBGCqjmqK/x9i455/TdbMgjmaw1PNvWKyDT8UVeYuVdjRzl1y86yHVGIh7w+O4yuEl
0USUxv8cBKPHL27QenJ3a2e+FVymPWJYWVco0HduXy8/qsXmtq1DGbCYg+egOJylYIO1ouUn6UMr
YiFbHEqOkqqT4BzUDRVTEV56ny6/VtPGnyQ9vRm9qF2C23DRv8ZrIMXNrsERmKi8s3/DaqbxNUuq
hwgfQHmaU8hgsVfdKd1PekTSngQlPzmiA+VOl27JMysnd2nMVqxCzUYc7GcGept4Fu582i2GZPSO
Qr3u+ER9hlMSyZ9cJPNutfG86AogIb0BhusfC04W9q0wixQF83fbF5PbZFgtNcsCd2BmadDEsM2N
fyAnQrN+CRRHJ13f3fIAkW42cAOO9mJWMAVGtzpitA0KZpJ0qp+YTfhbqyeDj+J0k6Y2lk9uyoDX
t+Grku3iR8JFUBt8dnyrFdMmR8Py7NHmucaIJrbYuMdglT/Ukbmv/+Y8U8B6aQ8Jr1X96n9rIVIG
69+4H/OMD5n8ZIML6bs1+y/5TEZkxv0R7fWMFC7Kl4IpKzeHdeDwrcvyDyXVWvVUP6/s9ryWdvSl
xBr+/5VjUuaUNPgY1o18MdS8qM89Np2m5pUi9+ucPIaVl6EilOI1vbRRkSqgR4YDue/cGG0o1A++
hxgdj0Z10pl2p3hZdJD6v9LKmAW+Rcu+RxUdVPngsZPMmlx95zXwCqEZU96wg7FI1DhuIt6KNhX+
+rdnUIoV5DeUhWkCqrlPKyBgn95N2qCuCJEew/h2eg922xJYJtJDYDIuLHMWTkCx9MQk7HJmTQIc
Q4MLsdlIa505lCugpIw3v/LgNE2P3GD7kZyNhbOGnvLKipbnp0xx7g2g1Vr+kmjdfrGCzhZsEI+8
Do6cUDD1mAvY0+7spW/kHpkruZolOpPkni0v28XCBOnHmzZnWVsF5jk4Yv1iRrq71Tpu1tOT1HeX
J4JOUI1x2SF/Pq0MWXXcNZKsCIxxtw5glPR06GhUhmIZDzeOt4g/vUNEb6WwF5o7Y5tN2h+YVA70
RtiiREj2cIeCI9G8afeaIJ2ofDYRO+Ww9T1FQQfug9mNDarBzBt6SOIqV6YjVHhvem3fWGRRl4ce
680N9qz2yF18yGtQ5YqW3SJGsJp/Hmd+XAOucvtmlLSt/hynk/hqm2b6ekvvaFknD8ZJ+MIz306C
wgY6adwgaEkyu8QUIASYwWw1PsMA+HfjGjybOF6Drgqdfbnw9/e7ANTIuCRXpPTcdH7MG5meDTx7
+VKZ7jik6Et6hvC0RSHYH4BdeHERL+k5pbRdTpkLckmjN3QPlv9P3gXPeGjF11hjWwM3ayDOG+hD
1y+dmAXOpVEn+6HXqjFpTPbKHA9+rZ8md+FlNjm3P22zGAbzR8MJcMqwUPhNa1oO/MAAnszWsEC0
yfbhvRQyZJ4wkQcb7RjkG8Y2OVbdfg/Dbay3p86uaYLC5py4q5ZuWxR+Sy91IzOyWRjx/mgiJik9
Rka8HWrrUQThJxh8RAknBo4RPIpGU0XjJ0GGTSUV4T/TNnMKl0sR1eMyyYPUKa3NBCpXbadJdnUq
vlgvCxME4vj99yH1UbLQta+5/6aG/jHZUkmghlobawoS+nj4vpJ/DI3bv+5bAme7CDFgFuyClAia
DosXxqlWpdkucYQu2gAS+ohC4HBoIuOMWuWShz+bWX8T/seTFZ7x2/fEQ6Kful7J5/6gERjuEtOC
45YbDjdrKuZ+BNZKZnh5w6FEO6Dq4X2PxjFcSrKBWGwcHNIA1M1F/QkmUZxAorW6D2sWKJAyfk5z
rkSj05s7oNFlD+2hJb0SFQGuE3Mh048iVFmkiXAIJBqWYUVzQBdRhNfS+NXTvcUxKTHefgGQ+XNS
53JDBHBm4dVCrFSQ5nHE50eMtYiZBiq4kCBFviUPYuxC7wHSpU/PI96kABdN130hyC14N1OkU4Ik
MFG6FBdast6Sdb2XbO4JOuiOT/VJCndrQgDOPG540diz1uyuTCXv7ESvq8uixY42TP2jSvp858ID
l4gAGP/bfh19cAQmX633gNzmC87L85ZhBNoSzMrICOO4dF1kNNELJaOfVicHJkrpSXXjlUHfrPuM
xDRSMzrNuwNwjil1Xs9LsiwDaO1fpv43xybsrBjz1IT19Lbs+MMmsAjICiefA1+s7B8V3MmYGotL
zhhFgqJ7HN95iqNYxjaY2KiRpPjWRL56XYSDPlMMQwvzqsluGol6SPUpUND9yZq94rRdTuUTGLLq
Z+o0QNLjijuZ3O2YxYe4PuOvJqWi/iPtDpdKrlAiBszXWLOB92qMYnwDyIH/hJL45i8jXIbGMhmd
fjgWBaFXWmQOMsxCMzf3YlMcck2BRl+boX1Y2njzLEwgNs+gmdNVgy8SuAMLfFrY3ZHfAm3nJ7Ov
VajS2Tgvi5OhA3xJnEqp38wpvVkYOy1KrUAz+y7fKIs20oUM+ZBDji7Rhecnj6YspNY+bzgK17OZ
ZRG6PhZxCgErm8C+h9kC0VNvyIHRQVJM4jy0GwbaYHt65kr9yrfr5iSoGm3Rgs9D95fIbSFWyDyi
Yqy06euq5PBLjCg+iAtLnFeJryLpKcprPopoKOJqGubjrv3mYI6nLFe19BQOxkm3weaFpPu9uFoS
LlDNBcc4M+LuUAxf+cYYUko5vFv68g6/c/+uXwfbneQCdrRuUPKvqLamZJ0wOuzixR7tp6ipKTqX
WcnPBonxzPhSiGoo1vWUnWs27Kz3ORJ6/wjRlAEalIkYJxMcaUgtkZ5NP80FnvMGFQN6rLFl9eUb
yc114dzNq3OuUtMuAma5jVcVw/YzWT5FMSvwk4oJiKMzuKHP6kSFgH0zKk+3gioQE1EFutal8H/V
OtiFbac4E32GN+r5+Tnr9qZdhbGNcITsEBIBPtPuC8ttm0xS3G13BvoZn0jpQJ9yzZW+9EJG4TeQ
jlBy5bn/5o3GSbtImCw/x06bkOLJJOChQddmz1xS4G++Zm9lx3gNjHKLrlTkckTesWsBJEVHWshA
G162dn87fldhs5WfwrML9cdcup77Jdg5Nq/yirgs1z780v2QCZSEqE0QwET+H05SwNC8mQjAFEry
ggwRN/5sJK6rOErnNVAYLJQd7Q9xZDfgjkXGmKCBL7CPraaReIUFnZiH69Q2OK9+4K6VgywB66FB
fAVR3nOSV710xFOEky2Y7VvrcziaMgVDJv+AbzcGiChqy2LiuTRmRAR0e7gNhksQXdhEHZ9YFozY
U0ANLOMlJHt/WagtbRQzBEtvc30TZz69sHlI5DS3JA6yBlWbWo+pauUerNeiYCqOYbVcSAMI7xWV
OKi4akXVpXgkIky3As4SYsUc6f4riYPWubPTPWVPbDn2uek6EkRYyOA8NqYf29IFFanBqWQOMYUo
XfnpHfzHXko7Ay55kP33C/I0hzJnqRJOenk1dX3UIux6cC+H1uPF15JJUon5rpAcwwtGUrb2yyv5
k35XkadvvJr3FJcwNnQlB7Bw3+J+PQY34y3+wF8B0HDm5z1xEVkc/gA8du/LldtOsapVoBYaDTzP
+I+BdDVUNqduK82OjEFAZKDBzTHqFJr8VOasiSlejix8FG6Yi5qKOK61XIskBY+NA9A2z+awRz12
b+YJ3osAA6MWtJQ2dQ0phCvxuX/n1jrEstWJ4JbhAasdBcgPkEpXSuG55jWK85Xt8jsUisAKmLDC
RPC9tjMLi6kuZ1jNGyc72rxWoroFFBvlDiAFsC3RkPFPpjxh+kKrVdcRODSTdHWWHbDECQJGbQ6l
mNUOlAySscatfBDlP6ggdb4Fs4Mp9+e9EIth8+H+0dhxIstxzOubOYQ4mk3/XlEbp2wqClTD87HR
3hCcWJg6WcMUVIhb5dVV37bVzQrqWk1TIxJ82OjA6YctiZwz6MhtDwxUztT7vXbK4nQwdhafjI3q
vssD/NmKtdwhH8rVZUMZqp2XaE9aWmMdcDB6phlVUyIj6GujYuAzDb699HGMG6d4Y5l7vQTFXbc1
Bjhz0BWMXhcqFiD4i9JnM1zWLo/pXZGc1xe+uQxMEJw7d6EuYbOQUFDe6Sp88gUF4MBaGXpuzBRD
lN4EdtwHTvu4LWkmQ8eWUT0SJxIZnTxzN6IaAyvc7zmxw8pcv0rwXGZNs2Oxwx2WAGmk70pM7fMU
OaYP4dUqOp6c5V00K3ulwevbAhS8ZRupSgcPVT5D4o1Gv1OlKpEpcBcL0I97PNs6BzpeMTz8fZKw
nkUmIA+uE4+z/q6zGE+QNYI+6Kwbunkd8xB33jD/XiI4AJb8XohLQ7949j2wCza6wDvTUW+6JhyO
d5SR0FLgdy6Cmk9TsbDBHEqVbV8JM7/U9Fdp3wBdJsVWASNeQ5gPWQjJjnjC+kcS1AKQGyJKkuPv
Mgjs2u09GRcp0OHvXZUr/VFbhI15bO1tND+L7TAmZcOB43LYLljEUj/B7zBbS8IcNmrlfZbIeJyy
qtHJIEKEoavJAh1bbOgRRbOr4+yBdlUVedEfdzW5GbnW2ncn+6MQlNWulHu1M5XkUSl0eJ/Lb8Sy
5WZVm/3syMqBjKF3gckyInaWF3E9DSDMWRJfGk0tt+uxCsqBb5sfOcE2jXgmf774dWG6mhdYeA8B
kvPUYvDw7kNVqoWI17CcjeO3gWGnXWtgWk58zqZrGWvvNWOAZyCIZlx+cF6Z9QZnIFJWDGQMKiRe
R/JXX+iQBMPD4bDCBbzYwIGL9JgSQtY7bnLmsSdUbLZ7PxANahqemrFkXBLQroSEPnbDVbDpao7Y
8jotMvsSZuKOLwM/vmSTP+YIBT4koek9sKuPfNZFFEdc6RHnxlcSWWVg55ipG4lf67EDHTnbzuYw
CVM5FZXmN7MFNHR7MsaTD5EnvLRrX1XVxRoQ/GrrHjOa2+j1nct6WM6G1L+baVP6deDxmrPGRhY4
yNi99MRLI6qXn3omyWDIq/w3fkUPwQRTE5y/2cqj/6tLpn9TbIrHvPDRoOn8bwa2HqM5XuwZBueQ
2iqmNX9I1fS3qbfBQiLTWDBxOHR2cLNJfLMLFzBwGVf10oDDb+omczNV90fnfZFgB3757r2gxBhL
5fR04E6ya7/wyUUwYQvBrTZQEv8cjWN4/5SG502OjalOvyn3sdaO75klXBnod6j7MrVgv8Nu6+Ge
nueID2O94UURV5v+EoX+IIHlojD+2bGIZs10+qp7jsQiIfExrotiYrMUF3TpGdSoEcIVGV4S3eHd
yIAMNjhSFIk4l7NqgDHz1q4rDB5i+Ed6dDfqUGdZTbDYRNRl1GmOY3PAE5uK378ZEzFFBzGWWW91
8bYHH2QVXaW7m/wEgkUmKNLR1AFLNBXpBXcjZE+YOjXTLEOi2971OA3tuMYYHNdPIBmuxMJ4SAq3
1fJlyCboME6AOZimNgFBXR7L/cQvLw5kgU3cYM2Wxcm9ksqu0c5ghemEC+Au3H8hWMm+933Ss4ZY
ulbaXMNvsAjrQ7QnKeSnxg+xP/JuhqdPS1r1G4Qqawm1YYWfS9EHKk3fxqugy0ejYhOo+vPwL7lo
6Kd4S8X9lDCeAPSbL7SXPyrD+sQyYIZPNJd1ZI4JxQVZ6LW0wqMTQGOE51B935omm7ed4tUiyEpC
y00Fh51zhWmgDHihgJ06+Fjisod6rqR+gu+ndcREqXQoSwj+y/vQd6SD+uCDyuKEIz/0yLs8h1Je
ftPKIRv4OBHHuFuaEtnbpDsI/+Bsu/yAE/pbuO3sMOsBP54OhrplYqkrGc+Ja5dVKHDzeCaQyjPU
V7hOtbGPm3lbYe4BcwY2EWTG/tYor70AncdBg0xToZACP6gsx8KBgVj4IE9SweZhkqRiDGk6xFVk
nFI8EKquYkxQZxHEK4b6tdMA/p4YCi3fdSd3hYC+FE/TEwj3KXfXch0sE/uvMTYlKzGtAGiAE5C8
ORotYP+drTT/ifd4uz8ZONYPyZWYDnwO9McCl2c9W+l2h8+Rfy6rUMW3GD6/g5Y5zXK9i4Yvn6fU
JGnpLvObrCxOXobl3Wcqipb8hZSfcFfTgCVlUCiYu38HGjhBrlB5Lc4U7xLWUYmwm9SG5dNLfJ72
k8Ilqt6zSQ6jp6U47s3ubxJw52DQoH/88Y3D6IBJkXO1m30kJr9tX/Lqfma5s2EAHQnAhJy1q/c7
4M2k/umfIMzuOCnhDWHnTG9gi4PG+rKmaJNhCgpj7tmK6Rip3FRyATlOjU5ZzDWByd0DtX3pspI/
d9ZrnPC10atbpr/OG9+OpdZimviF4bQXT0f5d1GUb9PVnZHtnk+iEY2p/nvN2fxbsZ2Phj/BRN50
QY0ici5zjQGNFFLC0QMv5nfw17q2YqM37zL6aZ8acAgqlP6sBLEMF6ant7VZyY85zgztpU4wbgPZ
nuTmoQxHClV+yVOAJ+zROS8+9j1VTRvYNkcWHJPm/eDbdflTP/y4L9YnK0spaUVBaEmpsr9qzPjg
nLmLX9Mva82wwFlYOh+mtZ4Ol4ncxi8zmbr6LJLP1J0E29A81ncXHLfQ5kRBkUkHAGqJv3ynrXGz
I1TK3cLWx0vNR4s3mk7AdD5rs7eWD20+qitXEgzqLc6oZSOIsiq6OpVjB5m967o8hrwtJ2fwjup+
Wwc0kJTM5kW9y4PSOXOJQDnGScQKaihoUYn+zy/wJwU61eqCrwek1FOeP4vYLrGVgqUPSKKn+8S6
Uon0zZHyqMDDa9J81HUhx+2yPMH4aCQD1t6bXId/4pnEyAsTi/P6UkHCM3hEl8KILwIybDPBYWcP
iW99Z1vR7DOIOOX/nMhSBK4ZAqitTH01iDxUX1tr7v3gFSXIJJELO+jm4HV3ETxyou2RzAs5bB3U
RbdukNTWpc9OVibjfixmug/iuZS9KxlPqrMOQ0IDcnawC7+os6ao9A6aqSekcIaqpNvkoMyj/asH
5bNnBH98VnCPBCASc9n647bnL5VEVODY10JCDXvUzg/dqwMgGPjcErGD8pAIIWHfMDucon49E35e
KUblDf4IGHWb0McpDBDkw92Ni53hkVUUN39m9wgRMAbQU7FbwHP2YyewA8FCn59VJyzxnKJTzsNm
kcSWZcjHbL9uWPUKOkt9ukdTKqx/ghciSQWXohPIu6qoQ54YKi0bR55QZzWl84VnBZDfk6kkk6Hn
WETO4F/6vqN5bJK8wv77RwhfHX7cbqqXZ2Mru0WaWHBX5Zad0+gQ56kGtId1+eMlWhNcmVxjxjDa
dwLDGvHRjtG+hHa/8oCMr88vsHRDFChDtKnouPsIZOj+MehDEFp2GeXdRXHvVGa8+uYAAHdMsugc
hZdXI4cL17S3xF0ftZzf8GehjqfqMcjqSrv0Vdmb1r5GpngqzO2XdU9Mntt9UaMe0AwtVwO7BDcy
IFxkozsI83MFr2xG27E49CEa/qHt2i5+XMdU7ZbAVxVMLaVJxxJGB6ej/B7Q2tV87/ntcF+VYfKv
uBQgiE6XVCRPfmEsdlFUgYrgxdZ4RrhvT94KUf3FXRMxRoHtePs0WgrMRYx2ApN2hs6PfezHLeQu
tS1O9cLtgKUKihw/fd8T7HD17qzmjvl34IZLMg3GBApriZxyr0glZGkXJMbKijqrYidi6z0uoeRb
nb66yEK/zxm3Gtu3sJ4AbuJX+9wupo6/LR9BKEVFJVZDd/0VcSakx8B2Kb++YyI25aAWHbAPQALu
htpXna4iS3aE+ag2ejg0LLypwjDtjv8MnHNkenCKMi+fTEzUhBqcjgY2p4FvDe8G7u4mt2Q/ThzF
TxJ4j7Lswhi+9wEAFkllTwpHOdy+M4SESuQBnacmheMA3bgkife2bcwDHXeSGwlsXv11LBT+bu6U
gBY9ukhDwgFzyBlKbuWfqwrqxYfOcKn+acJBp6Tc7Zgw2VuYZNggFlHYiA79/H7QPMtm3sDm/mrb
FN11TfFvK64T/6iUKOVTpS7pfMggdk7iRDLMYX4kcV2CuwZ9yUO6WaR9O+8G1cNG0LvVxA2g1gUp
HhrAFPpfFQbUHVDkQsFZEOXFBaARnpxiXTmbKU1rXZxdKfdVRHD/yGRiEceZ/6RXKpPKXqSof5Cd
xpvXM1smeG5GU0R7wTKLkawcwyKkEIQtXIIZJm9J+SzrQFRTCxRRCPjr9MdHAWo5LYjh0JQKqUKY
ThIVpGJHSD06NUDzkm6h/s1KAW2TrxC5+ps3b6jNdUBNLHRKAIGWYqmxPbqVGYwrZLcaETt2Q5Tu
nSxLh1GMZdupIsJd9Eqokjcl4YmUBbH2FSdN7ZLq56UYarwC8MkytpKx0PGuIcbjDzq0mVvT0uQX
yqmQYCKNfL14+N0/3pMKOxoQLYJXFxJUyb63suIuDynfVhP3BvdRaCoWaK1LSrab6dJ6w4G998kP
nrNZbHbDnzUboy19r6EEiSeRmL9z6VdnsRGr5q6Ll7hL8lZ0Jk1HSk23wPrPpT6vITq8+TCEQ2Re
Et93NU1Q8a/tb7UhS2yhWsyaW664XdUdkntlzsE7haDVXlrd6GhyFBvJ2W04G3u6crDrst0T2f2D
PpM4ZPd0nLYEIO8vfVuRkaNd2Xbp5kHf06nYdkS7a53ZUVmMZgpt/sS53qEjVIsaz09LYaQsY7R5
z56YS4Om3AwOaxFdPkbiwZNR10HGU4Aw/eBH8AJdT50aOzacP5rX9qgSU3hhJG6hgfWdgnQOqrFy
17pyNLRXXeUEv2Kzn4LU020QVEl9Re0mPSK6TL8gkJiZkswhRY2Lf1XyoLAQsmsT068wGI8DBVzh
l9BJgmqz1WIX2ealNQfR55qDsls5KP8I8AKjZ0ajl+Ao/BaBD+azKChDfElrs0hJNHCiiHmqVPb1
DMm//y+J7I9qyAKDPORS0e9zNyhaEUzA3jMxofWE3Jl+PgnPVh/nfbLVYl0onlDe5BRwn6o+oEOW
mwxsRQgnIQ91hYgILefDxF4GT34SQVaUp1KBtXzgu413PStru/4ZGc2zocyc+VV6UGKyBQUS5afF
UVuvg/qWPonixglmRcF9AR1NmjXElG9rVbZ2lzie4xy3AB4NOXmS8obsq5ucqcPGA1p0nLLplqYC
bPgcSp7/FkilH0RFlZ1HQn9pi7p58DyVYZ3JZrfDhB5boygYhPd+4ACBVZqsRzIMG+ib+N/Aglao
0O+J7hx8FiKru+bWiotxayAB8OX7JrNxBxC/GPbMoB8ucZSAPNDEwQJGZn9SxPS0zc+fSsvLMxhN
4D0fEXQk+mBTduMbJ/J3TpbVRiQuDole47hzTBEAOs9yzIBvbpFVZ5G5ZapZTbY4fYXgVWrl91Rg
hB9AjJ34YSXxnhssA+ouRB+k3ybUZgTQAEKAUWCx0AcKYiC64LbbIAXPAhqr2xGi1UFbl2ugkuB8
blHrpl6TW6smrajUHiUD4wBPIScyMHbCND01U59Xgu0zG5aWAagMOU3vbfML2F9to1QIXNNUj90X
TCPVb7uDfGB/1IxB+gvLp/kkAAM3C2ViIvaH27OejA/opWqODL5a5y/WEO53NnD//c+8+PO/qnVo
X101dZjz7406LhgIkIrGkKHS689aBHEPoaRz1+2QT1uz1Jyvwfs2mG1kkezv9smfNKk7hCmIuj92
WD2f4wipCMyY1PIhy3xpTj0rj4xmfdYuEFiZflPdFRPljpVgIG3zp/nTIeytbwP60Rdv2GazwldU
8KkDhKleNJS5OrfLDZMDVjq34+POU9DFLBXmXfFEDOACSLdDOg1jJ8+q/iYhNVvzTtF+GoSdd2C/
EwZBTOgcanNFZkUvGZ8JJ/N5/C1oC5AKlVZ8OxbdGDlxlVsSaFY1niZgA07j0H4EMYkE5cy1ez21
Wveeo2KszM5LcTSYgFZZbehdQtMJ0BK+0YxdrBnL9auS3/sGCRN0StrstJLBe8iSL8LuL9WBeZvW
57EXEyIW+Vi7Hb+OjCONO2ie+z5B4JgA9KSTfigJuApSqJl2XCUiBOuWfEHyhQfSIuDmi1Rn2Yl+
Jf0OFSCye27jOEZZHWK6LkFSHY2+8pgOl3v+Yn25gF+bz6Dr7q+JsfW4VufyegKEr/xUHxisDUd8
JoSN8W/6HUPDvuoeG3loA3SyUcD1kYwbRBpOvJB2rWg9O4GZ5Aabnu+JUmpksXSF1ZxmxoGMrX/J
5mhaSWQy4ylyoGq3oUEnXPKoHhg3u4d6YQ5JDgecwjSOeijbUU1+L1ngYb+EO9EJQA1mN3o+sucf
s9qJIfUJd1Rrxj/LGbIlK7v7JhiqIEdx4j5cSLVrrhheRa1OISiMiaSpQIhHN6c0pAETnocQe5EY
0bCEWR0XtKLOKWUpGZL11OBsyM2FqTY4gqxfzABrADGfzkGrUycNlQTvtZxCGzZJXXRbttykVcDV
S8nPjkQTCl5rqwOr5Hvq0GWVYhcihLY6AlzQ7mjfPGyKWhc8AJBhtqAKIsSCxtutnDr5uXNGKAy1
NfIMJe3AlL4xmBJDsm1OXZ12PScPe9ZD6eArgSbM50+wstHm7aM0lP1cEErlllq6FN29DqbbYQiv
fwT3muXElSfzyZI/owHMK09LL/PsgyMf/NiqTz6BpPL8Vzjo40i/6rBpq3ErbvtXBW4Kj5TzJfC4
b35KP5DsBgC18wFzFj1isO6UHzYKg5X52I/LHxzV7Ui0bvIRHU1yfCL4KpYh5Zn+ViviNaU+slXz
GiyyLZrDofLNtEBoyA7qUqGpzivQAhkg3IwxTdqFvxYEtiWpSITjMYVcW92EHTSX0J6wau6AkONy
pyUyL0Efg9ueNkJKWFUMH6dM4K/bZSc0oPNYgjJq7K3BuVQDkniyFhkVrC2vVo/QWF9QtlFleFci
kqiKCPP8CcMEW2ibVgbxBdXiuXP649neu9elmjZmahfSmdXhSnJmoyIEdOvJylG+2MUNzohswXgh
eJiYlfbNeJaHhUHxUUXEUBkXxKSk+zvupBIN1gHpC2R1sFBNOb/SIJQGSllCKN36XCQ1Cv+2it7v
aRSt/2GO3Lyho28Jk0+5JS8Ph2MqOlTPEhMAarzAqoAOZfdd9XdO91RfQTHw9Ae1l1zjLIglNYgq
+23+cUqN6WuPsaJsuyDtuwT9Bqr1lER2PEvg5cHBtafCgFVbayHyi1Z1wKWVFVkOkvJDyGfFDpMY
NDvxIxShoPL33elzsh8bqvfO745IOsYu8xmLfC+Kzyj3aPV1j3xzQXhiC1hZUs6KzFR87pD6+BFA
TDJDxKmXmHCSwN6GiS6+eWKpFvsojg6xlT2DXgCjIHpKYDs2aLhX6IyFIsmEzHuzMsxXU8BUeovH
G4d2CWKswlLMmy0emJyTeLqY96oMFJMD8BxhVxSRBFzSARWnTZbG4OzXM7PLSmrCaXQPeLmW2YzV
gRj63SyaNz1dMqDzrJc4+kSNStNKLNNVIsW6HpLu3RyXLVGOjmR/QWSl67gTaO8jIP6BmkEtMny4
LY6gu3g2DixlDZb7Q3srcqqvYldJF9+pZIhg5lpcjz6TYB/At/zGzewsTdSI9uzOOeMF+5dGjayZ
1I2sUY6dZU6Pt+EqcPYu+rap22AjJ1Q1mrMYLAMh51wDfmkosuTh8WFRafh7iAahUPpXGhhRwOZp
Cnl+tDlFygUU3l+S75b0aLJjZmLVism3JIG7gSqNK9iM8JRxkXTYljCbjUsMNRW+RDayiBaUChu3
wsVGgyNekMvX4iv62bJX8BLqsi4OYXf6ZyxGGd2Tn1EjsTEwvENRTHsoTcsTAoMiZYjOJ5wqAOHm
JZS+itaSOG9MJ03SOkCQJudebYT+RfNS84qquk7EfhvUgkLfJXSy8N5m76biVj7qCRlr8FpOOIoL
lwvIjwrMvBxnMKTJsXHiYq5j7cL/kroI4YoOhdbhY4F9BhIefvbjhJ3Ll5kUKzqn/0SU9ps13tV9
DPOMYFPv9jpYwdUsTgQ0DSQg5OuEu43Mni+0wlrK7L3G1gOzu5vj04CLLcfTl11Q/eWO/gA5ADXp
5g/9+6ZJQXCzM/uU7Gk8bF7Cn1omE4YkNPLpYt0zkT7CMZPdVvZiS2erhwfkw3aTFSlnVTJJ/rHN
pzDx1sfS9r6lSPUKcDzouwUiindUlLbDVIpFljfBe2WN6H7+/D+OTW5mTMkwjtKN4B+bpFWPowPe
/Qi+iBW5fl78GWTfyJKGblhTEQABlatwb3mKg4/VsY0UaOJ/tqs7uanc65T/rM4tMFX4ot8u4Mou
NnPwwFxTiL/woGn4HPf1SgIKGSYAe8Xh8kQYhDdwwqSemmdPvyEAOjwUAnIsI9On7EDi4eklnCF+
zhX3bR0+8tgyR73SE0dwI+Awrm5z+2ebWkmd+51fsBMo3uKkl6Rl+oAHOUmfwCMK2vBP6lj9JK9B
w+GOaxYO+4Ovh214CPTXLZUYSgSLikKZwqnGhNCnYHS0fdZIvViu0l2rLGTN7lZJFrRru52oE//7
MK8iLyNydGFWbKYk6ZKf7Khd9zHS+OGM/jLKpS/hG/YGryh+OGrtyepM/gtFAdu8d5LSzOzautr+
Hvo+p1wtt47i7hMre/QII2ihyR+Lhw5nZgjgdomAZPbBTio8rw8U8DDoen4ydC3LbxEF5oQkrGhT
pq3XqjYj0QMen2tdyv+QFBEbq6Zdv7spkhYV376bBBHTnu/5x96NL3KnhUn7TOSIrtj5WFq7zyEg
t30nb70AP/8hwXk2nCetUm/4wV1TK29XHdjgAbwTCH1yllIMkk9iH2mfbkAKv33QWS4glssTZ1lc
tzShi7u1vw6y98375gzTWH/yNyQNPoAJ2AEndgJH7YTvomXt4J8ImmWQ03K2b1gkK0XwA/gGpIEg
B4ZlmEv6Ix7QmRt6hoAsNsdozsUYfrp6yEcl4Tuz8FJau4mXFPsklodZrV/C14QCUkxVyv8V3J9v
DLLSAzxQRvrVByDNU3Vhp9oSCjuGs4Q7T0aRLUilm1s4Vixkcbmu++vfkNuFmeJCNv0ma23a27v5
M70aez7MNEHZJ6+nKzxwpwdviLF7bCKwB/MVmB6hShsbNkjB22dzLr7Xw80/MlXmoPIDw/PygVW7
83ymgYJKoVyEr0mFkoOnoQmJBzctPue+oIh3E5RR63pECQbBIGH/qKnJUVoBmd/TLDzns2tRmKI0
PIixsfjh0hoApTW2tBLrbmybKMUO2vj9smSfUmx8Bl/eZiP/C73ebaJaoTDhRjb+l3h/dvsb3FCP
ixGYXr44n2Msqsa17C/X8aFks5M+EMQLIfGnGrOvTcFmWmktD2S+DW1fa3aDRAk7mJjghJhaos2s
y1ds/s/2hd/AIXrmteRrhfPlFfY4MpZOdTjnkCKzA7DlJVIW/d0q+/qEr8WBq8wL1Gj6kZOShawM
9OTO/LIMD2IKjiPspjLDdn+C8mJsSjH1hS+Ftx1VZgJYujTQ0QIpt3m9pYBe6ub79PGP6wyFLHF1
xAyxPfozdwU+1w9GLL5c8rXIPVzJ41hGY2C9vJ+Mxr0deBZNMf0lArs1+eAJ+k67PexZCEYyUOpW
f81jzDGeuv/4kMieWYaCnw4YEWfq4mrdoj+VusHov+0H5uI8LrfMExM0OiQgwAXKFUlqBZSe3Ep+
VJdsBQAsrVo9BRf7l5DfBT8YjYPv2dyNV14Vi6yavdqBeZSu84K2qjSu2DVA6ZekRFLGJR+kqZtQ
9WbnsxretMOyFU+P4btKAz84lQK//6OgusgjiitTcSfGh4byh4sWzg+L/ExD/NAPFpFwYoXWZi/T
sVo4n1aMnkXfGmd1xy1OHmnj+CLWCQXyEKDinq7vMCY0TMGxdf/4R9QVQLRIKDxPN8j3EWLuyQ8T
dOYtrhDnZ8NWvM0TxoB0NO+HlkreIJZk5rOQMSWX75r8akilq9BMV0M4rssB438ZoB2JrIhh86Aq
fAbSLdNacWW2DAQCSG9YMNdZ7W4+Ly5KbBSBwGv8UehxyggtbNolcNZ8/6KNXUgl2eXwSCicmmcN
OP3c6K7XI2Bwoy9eSmlIW8PdAlnZAsa+EiUuphgx2yMUrrFGsw5ZxxvSoI33M6GcTzyWjr57F2Cp
mSh3D2qpT2L4xPTRiuFpGjWmZDj7NLREERgeCfKigHIYyneE0P3A6VmNboiSBl+n4QJFmeoN7GIw
+G4AYVuXmrUnh4vlJ7/9A93jtAwCDTxaMgJxUw7uB/nmgnUbYIpfMs7C5Z9GlYk55jJW8HFhihJ3
DY1BlwhIUqvDjm88fuOTgXZ/mJvsjIgCKKmuVN2ZrpNO38u27/NubJLYwFJmwz1/vNvFIpzgNHFC
un7otxfa+S3rMp4PBMIYtWj4ZSEmvhnlbIqO1hZraKBFTMosdS81LDSAqdmRUxLJVUoWCp1GdjLq
Lyx3bu9GrwYMFtwyowou+8/Iu/HXVJk90NiiiZwKF0v73MaOfkTYUdoaK44vgLTxFtZHqDS6fn+A
Nkw6O+21HPAxz2Epv6aL3Lja0uoV+dE98UeiRzA3AL2gMbZ3bbZomS7aL/upsK8McLwT6HHM5bYy
0DkjI2iu4IIWfVAjEnSbhmqv5l86QQ6gvOM5KUY2HQh/X93js9g98UNn5hDot5HCihNpeot22aS5
Dl/pXeKK6furlTclGTp/qnzfZryZ9pvo1e3nxjHe2UJiQy3TthFQloiB2DVRLZCoGHbxspNzIhR6
onVOkaItfPliRW+tiu+JO0j6iD+usSIhWGUjCHzTKsITICxftbCh4OaBpRNnhQ5dV0NjUp0CPquD
Dj034PQ4ltGH/n2V7Qi7adOCX57LaucyVsKmlfrXHR4le3LQ2TydN8J88BOcXDgM5pUXecxfigGt
zUhmrQsORgAOeMtiNyIvA71GW/cZz3b3jsU6nKjlKtLnvag3t4nq2c3fMQNSvH14Um69fQNHP3TG
EDblEOr5ZB8mO9FEBZTmZ2ZRPw1v8LR/ThOM/6aN1f0ckibNCtJKcEH+F+IaxXSfkReF9QDanlam
zI/++0c+YkMemneocjYbiGGu3YvU+nLgoOPVie7xDnPiu9Mr1mu4onHEYi+sYaEJ3BBAToElMEoQ
Qy684FlyYJe2ESNTB0ZYBJM+Y4jcWQoH5RPiWqwWjlBG8qoVCLLnCbsXRGKOOMNFxgY8AeKLjK0b
VGgs4Rxkvu0Fs7+c7ZOzGYOJJD3uJy8M77Fu6dQHM0I//4zuUyl1UZGukdxJ4sVuSqS6Wes4Nt8u
RB3Edoa1+q2p78rnq/UkrP0F+IKHp+6/tHyHh42K3mNFclhF4y9O4C4fb0zbCCCwVR0mYbEk4Zy/
gYT0W0Me/3eoNu27Li0OJ2gDyhp4WovnXLoipJs6Dm4BwoFyY9mmX9SMTCz301FgVsJ74pdMLodR
kWJ/vupxWJKojAp3C5EZulZRzmUZHtJUYD/I4oyEMVexcL4LNOz003vn+AK7zHBwpIgcA4VyUT99
KBIY/sI8qtxCI9H8gObVHJDjRcJ/3+LSuT3aur3dxLmWJmdUO19mk5dyC5vK9/aESVsFjQWi86sa
PXpbcyQuQGt/UJWA0Au+rEt4CiyzGhNGsOWm011glmvcFshvzEUCMN4pvIFNXqSG9gnUHShuW3xA
21QiN5nV3I1CRu6HVXJOlX8lZTYqiCwNc9CCfWitcLP140gqKbkv5/aiEz0PW4cb+WHLV/DrjUud
rSIQ/+/aQZkF1uA+yvp+C4ggfTlv+CqPdfl6qLdWS24FhH4OwrFEmd0sg2dW2IpLfyhobEaRzVB9
7Pwv/aUKZYNhPcF11GFBNKucp6ja9RZAiDMYULHNOxJ0wvh2qcKZR2ZQrgvQ36iOXu+unmqwfFvP
cSJjK8ch/Mj/5Wljdy6bD0ifw1fu/MnaYN5HQ5ug1jRFE/ERvVZln5b7HzGwOuXv4tlnWP8pzQfS
UE5qnhTlQ0UCUN8U+OWbVZZmH/8r5tU7dd021bA/RelF93P7FIkD0kZ4g033h0hnwGk140eJT3E3
Dn3Cz8FMtRn/9vRrZa7exQj0kKVYdYB92VyXfjEMJgHCuAyETGKWPDzUO/6z/hPa4ho+ZoTBdUtd
PZcmR938wqIe0ucE8a4x0zSAYnhMVEC143gN1AknYJkTXxh3+jBbHdDTmNeMtmolCT2faMQEdU0L
Vp00LxuNfoP/lAa1j1MsgQnVouH9dLT9iLjIMUy/TSceIb72w1G1481WXPWIiIw0nmvYk3f8Hqkw
W3daUuh2ck6x4vrz1ODt4Bl1eKhxiaCi6cwdXBBX7tykyf22GJxbYQI2nT8UF+ZautCG1h7s0puZ
sq6EdEb2+oaxwggZCwdyX3zNlxgwBPXtJ8jRPrbTbhtmSOmcDF9rZz1dSihO/viFkfb71k7VMkA4
VsShj2XmPY9vnxkNiepAOi7qIEGFN2BpJCmFwmI7ZGhKafDnj0iNuKBC948PGSIsnefQqlqJvL36
C4tZ5eGj4ADI3C3dzVqW5DVI62iKMIw6qeQsfdhJY1E5XgWFwGekk0H6sV3ydUTKxVkmntncR06M
KuoXZojpa0sDyHvRzLFauHwOsOR5/j1u7GmrxeGk23Pn9D8rmvxvks/HTKo005Ct/ORNvy5XXpzh
WTWdoGlongGEqKYWDYSj9yD4+9WWLGQcHMPploRET8O0Bq0LshnUF37+7iCangs0Z7VG5FJtSA/6
PfHtCgmkUDlVZnda/SJR2uf1AIdFuZNnsoAVIVp/d2yqmAPpWoamu8r0Ma3Qp4JAy3atp4jN+Eeq
MB+prIRA5D+WSFduDcNIk2bBl7fTyZtHEkEablvucO4Q5IEnOdVuOhz8bpwiM1cTAwwer/HD0OGJ
4I4mZ+Xt/POzoBFNpE2ez5MPCiufHYViyPaeFRMi3DVhGq0wVuNFYaN4NscLlu/Hgyh9Ho837grb
WZDfbmQHxsCTkYvpt1epsZGqYj4fsOI/164dgfcuGkLanlEojsGAs3l36N/aV4rHnHDx3k7sKdu2
vLeM5UR18+rTLzsk6MULgXQ3BFRIqBIOUMY6C7zQqcW4x19bvvr1mrNWm1Lqrg8vQbwnLsyT6ulr
k9X2xeKt+4QveVpX4fcT6PBzd9/h6U+GUW+GvGs7v3YkIMn5KweBnvaV2dZdX+karp6NqXQfmM7+
mOVIkjt+9LBCcbVccMkw5LnM8E4DFzUBBtMmJLv3z8VhPg6DtQat+eT5KHPLnrxOt/kIqX1FYGJw
KZtAxdm+43vHy7Z0UsyI5Nub40Lb/BLdH5E0bzZ89vQx+6NNI+SYIntwYlbKSPyAUQ72HUg72eMl
R2ZVVAk+vsdHMRm4dtziyEGnjDPrCyvlQdl19g2vRZDIbl3ZICztxrZxr5x+2RraeI7d8hypRQJR
wWncFnjlx3NOeRzyPRQWf5L3yAzIZIVWxhIazX0UXB+Mx3pM9lZQaZSppqVp0a++8qpM2if0j+oK
Vqe8z7l/1RL3APkd6iZ98CDG9Iu3aBY7tBgxBreSYdGplH/4lFdn1y/hVNGGz2rkVpreEqKqV40K
rqKu8zz9NFpzEDTDgcZrrfDxf49KVlLoYPBmlZuoPr0v4Xk360pZL4a3NeECciPxrVRMn8rn8E7k
O2/mkI+XDjC2JSxe0yQ70zPHICC7ti80Gd81MOmYF9k063gdLfACmsXxCFgbIdYCr49TCxX6/TAv
t/MOE0LwNner7nCjCiKk2n+bM2Puk3kJuo9Guw3UFO2Ui1GljLDr6cuj+L5a5TW5+xI9DxTmypEY
S1PfRym6qM4ugy1AidCLNNF8TR26xZmeRRZGU0Zte5AzeEkLZDWfHOH1bsDQwlmkaLS7OFHrxXnN
okCLJfhxWRPgBvskDcKw7c7NwgAJWspM8QUUZZofEPLDRGK53KqfkoVonQD+jhlSfumvPTp01EkY
MvaIBfIsHXv+Ow/3/H1LN08gTbH7y9DdfniwXJLU7tnyZ0SrFc/itEF8beGEazATAfXCdlHNP1Y+
xzLuYFyc3uHTYNbum0OQNzUC9gFWEfrbJP+DIsm7gzVigJWe+HIMHjVLBihMs4E/RFlz6WsJ1kCn
YRb0Z6eDJz+yvM2b0X02RoB5Pe1jqjBiMDdNVXxxn/S2uzAVVRVk5paWcOZl/OXEZNz4UQS50ea3
TX/x99qAQyu5fD+LKQRucTAKCEYABkYEohdN1tEY4+ulob6RZBydJwQA7Dp7X42IiiMZZ7rZgWkt
NCOsG4XcFy4y3E/Ssk7M+ttyi9OsNJDAW0l3sjIGsoGtWL9gOYcR+C3Mws6vb0DtPYF6i7RSVICy
mqoYV+8bW0Da+cKlvw4p1Y93THpZdbmj1sX98DJNRrWtwD001FJoI8pfsoPg3s5Z1PmmU9ApX+pH
J59QDC479yJWUImeJ5muQKVGhBEEU+6uUB/b3WEfM2yXLVYCTrntRm+NEzks6OVeQ89TeP1Lm5Gg
RYZJ7DFyKD7HpXZfkYh0mA//dGSWb6U6lvme64bFsesHunqxq4ZcA9NCoeN0SZ14/jLLEclwDjDP
DqSsnD23Bb2j31SbM6NE5VyrG4/LgsofVYuRpe9ZMZTSGxbcTVtwWjZqSWlPlgHOSjn2gRNY7qvD
yKGP6+a1PK85Rnj49WwFGalCr9TG4zGJ2vaYcdZm68LQLkC0sB8A+zq+otVmdHPgL94M/qzAuuXv
qY6JSsr95rtLhsji1mPSkiS6Isj0a6ryUcgyoWi/4a9haNhKIIOgu4M3vbFFHqPsIWDY4YF+K6f1
zqxOG+B2+fhGvWDAV5/HAObRb6vi2TRL2NyVthcTMJ3gf4twRs+t08O4ZX+oueS0AEbl9FHkb722
oVbEqUVlwjiHC7LJ2dRIB5qivkwomMxL0cXpob+kfEU/htjhyRxzOeu32nRAlvfLvELOlfz00i5+
QSyXJV4STBGzlBd/nxfUtNuquEJ0W9u/MO4G9T4jvPytdvcj8k9aq3ShfoJWzKkpqMnBBgihH8sU
BtRkWyyfxdXzixiiP+dlPoADWmK1Op4toB0iyw1dMVFpu2TtzjWTU1YXxJ8XspuwUmw9yem6Rtik
xnSoTENzZ2T5gSGVqOupQE8so5pBGtET9dDZFClQMz3CHj0e4keRs+LAqprreguCe53Lwrp1Q18c
OOSfd/W9NwwbNCRjSyB9Huj6b6P9lRbHgoTRsM9Ecg3jWRWoKhAoSqXoHn+O6GLah8RKite8W4wx
ygOzzGHDITXuB1kxRdPX82PKY+lLr6WnQxcEJtSELMGSTeJb6z164KnQRllPNsxvo8vGveX1ujhB
W3NR9vXL9C//XP070Ab2boJ5/wRYL84fmiWs7T9cifUej2/LHYeUlcw19E286knUrgrPic0fEyTU
SUmmu1FkxcUOnaDmyISoEXx9xYYUzl79pCgIVEDtINnZKAEjOiUqcF+N4zX4WVGw0RpXjld6/dd2
UZnyLDU7ER1UTRi/4QkTxLwUkMfCVL65NA3Ejjwu/tyUsuPlcxhjf59X8vUiv0by1KcQUnXLpWKx
Qit92JM4YGI2WZQH1CzMHaOws2AZLbaFhD4HWXV4iv5bl0Nuku/ugi2dj/R+bvAeYGaAey9gbln4
xozH0fUko+PZmf0RUx2o5xg05yT8tdcH3/HvyBK5AoU7PfiFvqW9hBTeXzYjQU7yfEHnlAIeDHLF
BRodmshuYD5sFEv3hslvrKxO6XXVR97xs8ry45eO/V/lnTXUU/23CJeelhh8I0GMlVSBoVVonMNo
nKNEuDTaEqCMl/5qy6BEQQUsj1DZ7E+K/WzmeF324i5y2krSlgczaBy5G6ftjnJqBdAlThUyH52Y
wRND7yYv6d3q4SAMxL+CBXg0cL7JbneqHh9OiKH6h8Vo8TqNCpCKwsGRJNMDo81HvZEomhIOLdpZ
HQE7HcmN8nhzNHkZN47q2VNeda60JeSUPBBs0t73/jCCnEL84y7kmCbW7LybDa4SCRvGRv71tppr
mVolNNt7cM6ZSyD7kXBFQAPfsDgZEGIemIK/YrSzw40T7uwvhlCpsPMvVSG+eIQkC6NHJwaplaEO
tSw79vGXkBG4OAzIU16cDzZJ5JL/k8pLjHnUsV7+GAly3CNZK2//pfuBeVXL4VzBFpe+Yrrvu41L
V2CYmgun9OAyCWtubajZPHNMnJWwj8pusWwxnci0d+P0sP5wkbeRI567g1mQjox+X1CmKz6z5y7j
/Wx9XLWeRnHofZO/KGZxVFdGrwfo83+gBhAwcUsqanO4eVu4inP71xsLdsSwIza/HZn8clMO+qph
1lk/M0ALYsARvL4KbHRPTn5cFw5iyPidM09Q7qGh+JApd1UlJPACf1dvhZao7npUZJNIcrVWmpEC
Rpj6j58JMl7zs14cA08HlaEcwI0k3Pd5v08hu1yEJEjPRImOsnPq7WsqtET2DS7uA0iG7SFZABdQ
3tJgfGmtH9OuMKwXZ2x7vYOxfikCc/Iw0HVZR3oPIuSX3gizEu/uf9e/Ry6GmYF8ppQs+9fFWQyz
oG/1jNzj/2xVfgkr/LNegGcNwcxLvzKkUGC2q+eT70Ct1cldx5ImODIPygz0jx1IKc9w/p/OT7Tw
lmyMPJVp5yDy9kHpUeH/tJ8b9+80lJfGbP/j+vve+65AcxJvy0NssPFfjK+UXYiChyTU4yXRegQi
RrQcE8wOqinNqshJ7dNTT2TVlEKygy2glt/F372l8s47hFInXs1JjNWQQmLA5XcUoP1YIichzGz6
PubSHLD7tnDClGioNoSclRbBPAWa6qpSsD+LDfGbPMZqmAxRgy/NanoevPZiKYcuPShWPgel0koM
/WB4WfFKhqjaLqV16QRUyhFFuYTAbxApwmZzPzbb3sPo6tjPMiWSFBLhdX2MaAOY20gv+Vat9SAR
oM40jxtY6mDmy81OrCFGwjDefsigNLDH0OUMEPt0Z6hxAzbwlG49ARjoIj3CEOklCbPHS/4q4RoK
mvlBwubDM1fFJ5Lwtn7x/y4V1lgE++Bv0NcMO2A3zwYoY0vpeSATLFkB7HI1XMdcfnBOqLHJi61Z
Hua63M+aOdy3rd1fmmGTu9PmkhY/xo9rVciB0Nq2yIw3dM3PqjvveiudalRGqTGLlND3ssBunYfT
vFyutcB2r8GoVo4U7G5E6LQABo/SSE6/W+LpwZA2m0AGQpta812uSUfqeseclJ+Dln19YMxhogFS
jeKVQwkCPl4l0l35xFdLmOvykS8g5ukITZ7S/GVLdvIfUfZFZ2Km4Iylzz3DYhkV9rqG98gNwqDy
z5HZhIgA+qKUzjHN4L1+PmDxEP+VLoQGbZbAq53Qqtj4aOj6PNYqJ70jxfTWOHWZ1TXPKjz6r0oU
elCdHO7Xo3a4/aGsLAAIO9tv3hNbiUJm3tBAuVJ4ycFCxqJmsmpiLjMFgBII8vxFLQocZwlrwU/X
qYHxBa1FKqoTmfBLqm582bM7SAgDTkENyVcb/qm/iaGX+8S577Q7HAB454cz+UU+TLf9R0ikYlRd
SGUYejhTqjpvX/qkzDFk5+JZLvGCAGiQcEJ+02LGgA+yp8lg8DFB4vNhgoQJYaHN1zje2f8nIFjX
6u2XEcR+JVVqvveBNgLOxcTw/qlGVGMtP92VGC4r8lhTJOHtTAVTCgiDhutWCCv/MLWbeVhUmkTS
pzCeBaiWBeQHgglqCWpqoBvSEXkFHB0woSWJUGVN7yp/91tFH+dpRD89Rt0dbGkDUpaS+iyKzqTs
XclT+JQgmysR8K2YmdfYyB1yqBp91Fd8yI2QzaubG/mnvWbqtAzXf6k6rl0/2h1gFrjdpF582xUO
hVmnVCQWflsCBVCcNFlBshL4dHegbhF5tXL0LqzjX9yrVIunusPyGN7wapjmvBaTZBfw4OB5Pglt
PtBHU+Tjg8h0zqNx7aNvejTLcZQcYx7VimeilKfyvKmxPapY/wJwzzEapHuvFylJmI0/w/leOwkc
ijWgP5nAoHPDgFk7WpRNwBkKoCsiQa+Y7l900ZylOsS4zQfii1gkxTzRMgmj1bpvqLrJGGTyDMvR
Y00hPEDtKWaf8GvtzF53Pa/404EpLZepTKLrsyhS0BkWR7055W7zKL/BW/ek+l6WFImdU07JLbff
dNQ4a30hII9wFcS1MFDBz9DgaK3HiZ6OVZK0I7pqhM0NYtIYT5o2r+eA2gk1V8ZpLp4aGv4BI223
LFHeCBLwRzdakibCoR8qeK2OE5dMER/4qLObEmXJYbp9+rfNqIl19DJQuLprn8QZj1S7YIURnPlV
fZh8Efa+o/MnaWQJN8KK91b6Hi+bP4nUEUHTeGGCwA06AdB0A84hiHZzICw0GMcct1oxhmnFS9ue
L7IZxM3eepSURFaz6mZ34WF2GTr9NooFgqkuF98kNtplxTfN40HW6M8R/oW0cR+Q6vrDbBdEQAi4
KbCf20QtKAApxDd6Elp0M7oiEn9g18Bn6qq344/fBfDulfQmohoVrw7mpLMgLd6NWNpcdsChdQBo
qwlysB6tf9Hz06cqvMtIZ5N7GtObeSiHec+jSAePndvBQWo85s6895yIP/1UrGBmbC9e3o1dGk+1
tA17q8cEonNsml76U59xggEYbeBXIBE8ScSmcX6xhFmb3PflieGGo3z7ymZuPCVBSSl5O+3O7gkV
4EZQo1eI0927RDotngCZaspY5AkZ8xMARYhxdNFhZJNdLif20Iv/PJeyCV23Pmmc0evlB8MbLzR3
XPMos3DlFprcd4j920ENJgZLrrY61IPn638Gj9fXpZwbYtChSZeNz1busPqjLVwDTx21Z2cwU/JW
h94NkuSdRaZY6R42zuJR/mv7Jy9y5CBia3PA/WSk+mDVuCf7cM2Pc6mkk1BRThVKbk0VcnFegGaT
BcX4rU20Mn2vuCHqGSH6ob0/eaxwVb7rXcB2PJKRGU+xF+dWlgSAEba/Rlg+0miQwN0nA6IIi/VE
99C3k8jI8zIw/FfioP3dj3m4JtlYMoEzT5XLn+nGsWPJiG8Zgz/jkOaYtybNFwLuD1K7XkMOy0n0
4uTPzznCZJbLwYcreL0MMNyHQVja3eImesb4V/j8cApKYG90UadFuDkJf8JkvpNSbrXnAN7LvKAn
6LEA4v3yOVqyW5M7qIObmgOYoARa1nMBjQjQ+KJO9+iWlChwbm8ZL6HIR6f4k7yTbx+TwveReVt7
dES/oOsHH8Hd76dUDaY8mEs2hKHjgTHGYE9Cvi91olkH5lsIGgYfGaDIaHWc4ymvAXMuTOoNZOdX
VcHlPvZ2tJUu5NGYOGYPLX1mgFdJTu/+oP5TilNfhkxVoT8l/6pRbZckL1M1oz8KUN3gRf81osRi
8UvU9JFzlG4mbWoq/QYPai3pLs51KSGJdXzFvq/0/3Ln67ctEclw1fo31/mbrCId/DDCbLz9RXeg
n/XJqOWF+dFdt4TKEld158HRZGHLoBf6sFPgwCnhJ+W0B1vUfToQkIbl8ScyqrAJN1Yez7zKKn4U
HNl0tVsaWZuj+cA3EMB4Dm987VspMLhyfi2rg57GqUW8l6IuVyIKefBQigo0eNYw4LgSy9LTQxeO
UzR9oMSk6cK/pAu+fRfWizvsYqg0N5lK+6sAalx/fRAh+fp07Ukd2FGvLJfDn/AXGA4AK3tdC34r
HOIvUSiZ17IGeZZmOzyyxgTDzh4MVavydGuLMETFT5hNSAEmeK44qIZtpVFQM6H0FZfVsUAiimYc
7VgkjwDTNnZGYmsxur9jjFOrmlAUYUZBZtkaMdO0E9J0n55IkkLubri04Fq7BcPLRogvl1vx/EzL
BdF8+NmHIz4ArbBqeceTylHVvTHBxP9phlthOQgf8IYHQKpe8bO0cXpLUCKge4xn/e1a+8ZYbeCY
stcAdZw4QjV3xFhxAKB6ZshEZi1V521XHGYT08co71LNHgbRY4diXK7z3pLC/yYQFd8v5exWLplo
zig+M7p8Os1QsuacseGIazoxSiAzARDvMetnubXOTFUmRmfY0kdEstk0q8Ogl6z/8FLm4mp4g3x2
/kIj4VeSbPArIQmt6lTBC28KXtdtpiFLhVgfbfEA1VrOtpGEWODCjpuJeLYWkFXdIDaQsKhAscNi
JiMHaZxEfLzC6hH5ks+Djsjphv3ggmInhUAxR9jhW7jWjLiNGyK2xDaBEtZ8n8ZYYEyzPgBi8Z1g
IsMd01MtnB+tAYgFWqaGQ9VUxrNdppzL+GJRHJ8Qmpw5jmc2Y/elnGHOhER0aqMEeAflu/DYwwUF
CmKhun4/HpIDgl3ZYYGPO8a8OC7RGtm042CKRWBp8euhEk+n/SUtW0ABlNnReRSFo3iEwZP6eXwp
I61JrYvl6HowIDb1PEWUJmrBzee6UryVmZacAwIv040pvV0/NDGfnOfdlW1Qloj9ArWt56yRPs52
tOkgFXVKfDf6dq02P6eGt15XbDGSaUJQlEz5hBzXOsaVTBvHmWUQd6EThu1v9t/jfMq+PymbL8sF
2oDk+IotR5sT1CkisHAiOmc+UIbX2PDRvt/HLTqiHELPvHg6w3PNs37ZszK3j/5YKXKnVcMWQQxn
CgTg0SMnb1ruhhhBBT+bebwY3g2YkMBEYcybDzm/wH5hnhE2+RmMcv5J93mLgX5gMsS+K8RWL1VS
yXlndj74uAb7pioZ4A2Qdbn+wmdQGNSPEGwso4GdjeeMdjg6xZsTyJBGfJyUZAMMxf+XVhiuQK87
MuWQFuG6pbN7DNlqZgIomk6H5LQf56poESXEtR0j/5MFlZ4VASvhoJJKeOu9fdhwrl/vqwmhLvN6
Xnn/7EdCgolkjUvjamiC3yNpsBYiWZgL/Qi2maCNpjugL9jwNPRhoI3f86up7Y0HEv/JUb9ggmqz
dcBofC2lq74PWC7qgeVhNoL9nlUm6FLVCaZa43+xvsMHyjtSxF5+82dgcAkK1v0yqMVUAIYhkO+I
mQZBsadIisTRiGotJF/C+WrdFIHIvvYrypktuz90vZOIbwWTeS2wHqvE3d8nvPSUFX3S7+KbJXdu
aHQi8xbKb/Fh/ofdA7wedY9qy+YITQNjeVrKWxv8C2Wxdv+XHqxdpzKRP5EzaZstxKp5RkP5JqAY
lSp0EDWNlRIaCVi18b9swB+xZtHtVjKJSUlEn60NJYEUphRtrEuBGNuZyjxowjlhRbT0eZ+qjylU
dxd0FghruPVYTBsqTj73SRlxAdYWMCGjZS+Sg8HbiiiyS+hTeVX0gs2rd/hC3014yBZl3butBn2W
IjFMny1JWtq1GGSw6zTnA3Dv6wGx9cUZ8DdbDOj2qchi6NArE8p4+evLYD80iL28C0MZ0FE3ybES
HTLAGvJt4frSH3XE84W+6kn+vNdoypSMkqB3qM/G5W7Hzjv2cucOeCWKPRqATlW9ToR0Bsw4I+6H
HxD4gmW0kql9TCulkIBHG9NDokZhLzWrUcD0OZ8Y1kpMh0NwyvrK8YYgo3ZPc2LnsXejIS7YyjIK
WBYS8UkQPi6phZcwMrEOfKE/qN/jUO42WAXG7KMz/LOcGnxYMRPgLxy9qmHHdhMUmCSPiazeiy4N
AZFijyOY/Xt9jBuY2SiEN66w1KNmFnPwpTyQUZaonw/O0jnrMHd9jlon2h20enxh22LbeBOJj8YE
MDhRJXkuob66zWTAxwG/kQwGS2kCsWUwPaassJ7ssF/v1qVWOcTEgVDBUqR7rAzBjBH+pkfQ4kH6
GEQz61zk2lddbiZlGYsSyP1TwJa9lTl+pWfupewevzDjmbsHpFo/nhAk3ZvkRGUulWqb/WAgkppQ
dkEAzlKaw4PBdCr2sEvybHQmT6gJ9NeFCHFuEe6L/OXOyeO/3Vprvwtf1kFNxlfj2T+b8fTD8eoT
0FXz5e8TtDQ4uHqthjFbcwqdg1lH8HPsKQYRlk0bsXWuNLRKYuCLkiyA7RQwIVkcphgyF6VCQSqs
npXn5xZg0fT0s4+fKifxkSTuYSoSL0XarSClaje2FGuuCHxkeGobPFec4D2rENEa75WC7kBQ5S/N
h5yobqYfJMUWdttUcliPzilLROjmkGVlB2zl3xplr7zGccpINSVoApU2im6KYIbNSCXf9Tt4LWJF
fQiMWPWAFuIQq/f++7FIt0lfuHpCN6PyAtcl55RlgMlzq6ALOICmq0m0HJEYOsuVklUnqk6SKXcf
P909D1Veeua6tlFIV4tyopTpdYN2MGt5arbrv2Ekwxj+tpr1HkhkgGXx0goWh7Sd19kV/IpctttR
UFRUFnF8E/m2ti2KKojCAK/StjVv/YqDuv7LyP428WZUcZelXz26J1kyuaVDzsSp6NseN6cr8v2l
fecHErRgbqafPlXdzCiBHWjE1Q2x+kb4E3zj2Ao+rnHmik0ARIkZRtA3Oh8Cqdj67H0ZJCQ6vwpi
BrHPOlE7d1w4JtaM4nKfYIvX0/x0FUXz1TnxO4vOgWcIy74a4Jr1ZXug1/aqB3Wli5ih/x6jMjum
j35E+wcUj/+Eo2wJ+6z6ZXEfH4HGBLlW7aUAkThJgu8nBwoyeCZcmXU0wAKx8gI7Lt0wXsI+1rfp
AzFaElpCIleqh++2u5ZBEZUf0Agkn3df8UhWZctSNCVsL5gt08k4Wu4KSbiM72eW/cQhwW0jh1vw
xxYdSk0Roqs4q2FhJ0lc52MMNeSQzwsjo7LmMqbj08i56E0TSCjjmqL8j10SJElFBSoNux8P4lQS
bdjwRse5TOAE2RdvO2BSkqWy1IiE3cRO5HRHD2qQAv2Ae5X2bXQz0QgSJ/Pxx+KeE/mg2mV0TyFZ
Y0KgGdUmUR1n14SZXJie+0GNZtKo1Jz7xQBdUpr5chaKxVoq2+AG+DtvSERgXr5UkJDKtO/0wzhH
O4aj4hAiy3kNBg40hB6KNxPvlyi7b336//9AMyC60i3KVXhZC5VLytTn4YCyP8elmSLMoVHGUdUS
NFFRyWsYVJqMh0MLBxQPKRFPlbfOMCEWIkz3ooMY+pCzrkEPENlGVeoEE/luN0Va4VP+J8dA/zgV
aqIdieKFCQfd132jFmg7gQTGGELxy8lXmXg4qYYFmxOOasAdGn3MfKPXN4a8CcHEN/7cXukHHJFT
wUnZzOkwMdsH/oadDQGBRa9rjHwwd/6EDkZ8TUXGi1dLBd2iV/8YXqrEAgX/WQCX9NNTG6x7cHDE
Vkbc0hjOvs6MTY5+MSTnHhX+T0IW/YjMQ+PTn0uu3IifQiIt4UsI5IdV2GiM8PUnsmYisi0GUSSa
5KIgjWP82LgovHZRyI0dr2gIeXBNv7yUVUUb2dji3sKp0LhC15v0Qm8+WTDRGrdh55N1bvwIE9fJ
WjauzygPXhJTwo8iyPuwnZ1GkH3xMdgdfKZ2h9HYpdPHSJ0A5uvi4KRMupk7SZQ2TC09w8Ovi5tw
pke9IbyrnBTlt9Ss51dQYNnLogfP2p/yzOwOD1q+9en7LW9DUGLim5P95dQb4Aul+NkHvcasYUJn
TN7v3+F61+4BpYEMQvp6GLpL1QoiujCq7jSizdbubOweb+5xXgnjB4MvP4WSN7lGvlGs/XkLbgcC
iWBVswhd/YpVuF3tBOlMOswx1v+D/cTLqvxSbkf2/zhc24us/l5eQavuYOC4pepq6+z8Erjo3gGu
f7rX4spiqp+yopj70HnWZLA6NQHk4oCgbawk4rPkkuiWIBKABuVFLOW8BaKhWF9Opoza+2bWGiNw
XHh4zDGiAwlWLV3iLwvvF7pwcXA7v7pfekJIZ4gITT8Z2frFMqVCQDlwPNqA6fj2znS5QMjy7Lky
x/oJ3UhGdn3ZyyGaC6qYPGAIhaZnpFV3v924k+TUDjBnpeSAwuWDp+0f6uvOlsP5Sa+2N3VCHBUu
vqwPlLEzXd0w+9gR0IKD6iFExhkGUIG8qZ9Cg0Tucdmfm4PTmumt+kysshvnnqsjnqzu0RL+rz84
gTuHJflRsOOx7MUas7uF+dHU9LW6oFM8uRppqLdo6QQPpUU1iGDM65A57LhYE2S06m1qC7MR1+79
PQ8O921uBg4egQtEc9dNZ66D6dYwZnJ5ZAjrpZTr71zwWmbcEkdP4pfGwUoDsDDaGLoZ5BQHYaxc
QCp+8sjrU6tVd7bBrFJ7O+IaqmEWe6UrVwcDdMbT8NNmN0gO6J4WNS+ux33d9+FgIrAqWLMp2Gqi
Vd3f7vgD0HDpbXmZMuqyRqZZduGPqIBd0zffhBNu79EXkwk+DIFVfvqs/I58mOuBs1O7R+ySmdKb
TMJmbpEHwMbODZIGVyjPKsIbrQWd7naUQQJ5p04Rjl6SlDKz0HoOjXCnX9dUQyE8q+CM+sQ3x6jg
eBMRp3z8qMbzupr7fhfkowm4cK2aeUt5v3ynzcKFfK6mttRYbApEBStt45m8yANGWWAnjiyvEL4M
TXmst3o/OAaokUMMCqVwJyuPJaUufdY2WVpji5DqKVQYmxAQr9yh92nvFTvxKh42h4ZK+9NSaUOg
MOYD5o/PRL65ZX2EfUD0RxofzCqrUR4ejZgsJzPMc834/5v+cN7yFWywETcJU0US2eDUbUi65QG9
dm0psfr5MA4ggIEo0K0oUSLksUW3FREVx40+UhaAsUhYsXPN0cRTiwr6cwekHUbQPddy7yKWaFOC
NWCByApSUV4t+69uF0SgMnowcmdyTuC5tf3A0EVCVAFO4BowlVbNlE57F2jMgRgigq1ahOFnoQuj
la/QqsnUgLITRRJ8TAibR3VYkOyJOsM+/1f/gQUUQZUNiAsa4+v9PwH/fWmxM+E2zzfqDuMivmwk
4M2JCVQ9qu9ETE3Rg6jIm5icVm/Bv3fVX4+RLnOVAnJRXelBVLfHCpDE/7LgEkchm7jjroraECuu
hALXJmkzfDgwewSUiGLgX73ISGA1TsfHT4VN+sKgT/nw1kYDhEv3a8qRTtwZ2169XMbgr8GNkB2R
SnJ1T3Ak8z8muXzHnMHr5niTFLguer5C3cwEVHsW7ilows84ZCFDSpkI/QbGM/bDSbqtC7LHCBzU
PO6Nl4w0A16LHtku0Y3Ti4r2WwSz13HdlXdbpcsJvWriTfcHW9zhyEe4uydQDCmHzkFxqStVlcc0
CkrVqlOdy/SyPZvdRb7WgiWZO+neOfCMNWIkfRLEEpfl3Sgqu2J2uXuTgCWAkFWPDzjBfBF2ymJ7
i3ZYfIrNXwB/LKUIFvcDkKoHZd2si79e2+s6itSzygqGo2ukYiy0JP0guRUBYJS/Ksk3tOXOLjXD
GATRcalv1bXaBeWrDtVN8cRp1vthJESd67VsLkxP6gefznUpvpIvls/hdoBrH0m4Bnp/3GL/K2fT
A9923i8wGpEFbKZkmD2umqZ9I3Bldbd2i64cuXnUKXP1gKyGggaX86xrl08dyuR+kNZabxGCEAiY
dyE09XACfkjExpTZ8AQ387XN4H6ya/gvV16RcxThhqQAin12P5itbC75UhA+ze1JI/OkV7OUaWZB
McS20T/wUv4mucZInsIDdAhlF9vakAKz0q3nboVJ8kIZJFHTf50bdLCqDgO+XHpgucUpCIknfgCI
WOqsAkMBTZu+HAFkCBd7jxzsNbz6YFRgVE4Sn9litcgjL1vxsMMH4tnK8WkZC44SMmL3WuqqQ+j5
WwW2nv/u7l7q5kiuanZe7chHu7ivlnacEUDejmpbfZ5Y608DtH5RtgwEuxK8DemIHY0lAaRCtu6n
psCFqWZWHzZcrsV+iWtznacPuHuMdTvzw2vmIb+MxdSOokZKK4UyzzHQfItGy89QhHH65w+UI0TQ
tc48TZw3p/H5Cq3r3CFqwrBgA+BWuUdzVV88qP0hbUBGmScyz+NfgWKMGPL2NpXpL697xC4c59zv
wMRFgcnmlR8+JuLZNJickXd+3p7OAnH+7I5LjYRjJNRQxteWed9F0tqM4qEfiuVr7ZWaf1n9evgL
VEmepV/BaDsc9CHyQE14PfWvHbVD1qzTphZ7y1oSIZvAZq1DrKEPwaJfyvnnVcKhJ/4PVBtpn7lQ
cl/kLufXC1VtVmhU+OEOO4B93pVpzb9aSIC7Q9Vbqm8hwbMqynpbMAGDEPk24V5s8iX2xM1Uha8k
XGl8DeMUhH8INTz8wa4wlPLifdol7490UKEoatEsXFr+QXGu/m19HRM862z+4f9orMb4kHaSb/1v
Pxvy7auruA0oy4YYr7iUjEwvHzfAxCWPG8pnsGyaVIvVO7K6c53MkQG/ATm0VxBcnt3gnr4QiA0b
LbEcJPVUv82SbUUkhG7w5qv2CAonN7dG/XEBO4Xj2CFSjD6bC0bGueNtKnjiEWIWoj9inTJlqzfY
Cm4G9PTNPf9xXH6+S8lwjSm73WwCp0fGnGHIZ+tid1QNjrxoejVUBMcNyPIc9MJdvNO4ck9Zla++
9QqoKRHFbrHh/x9/EtxRLrV4TYkM0vNOHoyq/u/R2uK7VGxApf9Zu2TesRhgoeaOl8CjMnI9H9A5
bAonFQbG5pZ3LA6Wqgfh+0fuqbmFJiC6Ji9v4bFwFPijXfwDML8QVPduKwThLcbCdAM0SW2I4hM7
lCv6BU8tYk2JBce29gKNoliPoyoUWtmKd56T7d17/tqxry2XhO7AiZAT32OUFc1MxCuETf8661A1
CtIu346xMpzvKHTxeR+7fEhL5/T/I3vWwtmMWMtofGZhtDZtmbgB5kDxhhru/4NWf5PSvazm2o0O
IbCJc9FmkNHRUHmEs67LUDbIvUL+cG1jtv+Z3jnLz3KW2QieamPhPwTXdfY7cTc/EeMPWfJTbLZ3
xyLfuADAiw12rBvZgRJ1Q49DL2i6HDJCl7tNzaA2UBuF9ztu2w15oZUYYHYd9LbjPq1fTTi2zqvL
y+rCAP6QyS6J+YoI9fihy+OQ9Xk+ij4AMWENxsPhLgN/36WIb2bGrYBvT1dKxR5B1VAeGLHboea1
V4kyVpbqpDh4PVOQhb8QK8IDOZUA8W4+W9RZULIep9QVx/ClJLPdlgMm/T4IKTCQwELnFnMjh0Xt
+GV/E9d4JryFdM1daED2Lno2J+eavNZ2vMQV3qf898lCGzpgBoXOQzErjud4dJqtahVkBABB0Ca5
DPot0MhbIuNpATo01ZbCCVjDmBJq2Z12HmGnrDm/BGVggMKp52WtLevTfNqBQKi1HG4bX8XjiE3W
gXSEQib43mg4KFmkB6RcljEDjySOuaguqxUYeKJ5IW7lix4ZHqCCRva6OLjS7JceyfOj97/6uthh
JrVa2AT+Iy+mXTsqdMynRPMfKNVlyeTPIgs81cwQ/BTbzCWZGlhJCaZidlcvHiyHml/FBGBlpDqC
AULVKHRA4cKmeTsW8elr7AG7Asi9WlsQ6F0kfTH49KoyvFHyzXeLLZDcidbypP7X7zYv39iDkOrm
RvP8LAeYcnT1CIEKcvj5869VqlQ028tu2enO2nv2Ho7yBT4cofLLw+CVuOalo9lhRqMEfzA8BMxM
lXuAnWvYxeHCYwkOtxtSfSSSKLUSUGArqDZG6bJ2vh4PfgVDnfc8jPI7Vn3XoNGSI2H9sabPDdso
3n36Hw4sgoZixqrM3v8QLj5Ra8oowzgIOun/kRLpFqmHYKRhjWijjP+OQqbohCfB6PWl+4VjsCKu
BVuMM1CPgr7Wa+QVZF7f4f0gI6ZeFew9z5dHdHx0VfEGYtu/qISRzL5x5Hbg1CO8BJ93+pbc3Rqv
p/evHaGUYbFY3GKu0G8yAFG5nzZrPJSNQiQbcti7q43ezADZBsSzkKsqPW46TDDMfYSsORgN87uF
XMOae6BV+CqBXgW6wahjHRsW+bAtY+y+NLMRIfAnOBxy9TiahogVeiKP7eHPDaPwltjjae5Qw64q
srPlWnNWK6fjof/Z9E8VCjRenlhr72qt4lrojHsTHWWoxj+elhAJwsYqHGjcB7uikngXNFP7TYPC
wmlboHv+vaC83N1zCFJsDN8X9IJqwGZ3Gc7Kc/vTmUDyBer4ZQyAK/yHpsNnYwckucOPxkXjOcGb
c226Lyr/5FLaTEKJaG5ZHJTB/Ys4HK3VFaRlq4sB3H6wdKmQUKBd2eIc4KhWN6u5PgyK9ZbDbhh7
gcvhveyh4Z4OH0jfIRv/I/b/tNMIY0wdmjvFRs4BNdVT+GYx31Lb87EZe9H+G1750SeC8mm4M0rG
+zd5hcYjmUEU0umOo9CFpKosTi5qTdRKNX2dmBAmOYcjuG+qfkyZHZVrtpws20UBrmCeHNuhRZeU
gMSRj824Wz7biQ6NvzWVQ8awT4cb+rRkcQD+TqrLto+r8fnusqf2zzyWhzzwZIy3/lS3PNwJmk1f
M5E2qTID8cHv5JuTqZCmzpbTW/g7d/PHp6rKFG4TZFbBaVkFhgYlkP4Kj3sqUYRE6SpuAHM9VDJE
b0aYEmtVR4K6IX9hj3PRBtT7aaNHRVEbndFA2+bMVPeYUUMHvhoDksPpcuLx9pX+Bsphxy2/UChm
bJu5YwEt8xwIpHJTqcyN9FdSV80bPIrudw7+wuqXkVmVnMk9wuLDpDXIqlZk6QxqjzLlHftkStGy
Sg9B1FW180D3Di5sSVSBI0dR/IqQS8dLLD2h+xChc/FUNdZ7g83kpj+qmmv+B9oqnuGsqCnfYORa
UUKaPEONLHeyMgWncFyCw7xNzPthqlQmG0y6+KrVufJwnVsmC0igacnGs7Q7WNhk3mLYRXMQ/RHF
GHzZ/G0hFUc8C3Ee6o+nFR/PRYBteCm4Qm3Wfvo5xLE0ITg6s57GyBomhYqaIHyQiDPtrvr3A6mH
trsOzFl7TtD68BcMPHMqjqmqt1yKL1SZO2uKylmBZZBpBnGYCS8P3iVVSG1ZkFedbhfQF9RqZeHZ
/jQrOFBQWOoTuRtrCu1QjyTWnIUzmw3Vb0uykrBzuuGwI5Xv1glipsjOmGY+1ZVQBaNXVuE2VqgU
YBX2csgOYgftFqaIwX2A3hIM6zfBduZgtS4K1T7WHHN62ZZ5TVPtONgWiljuiUe374Hrq1EQiQoU
CK1oUAKjYw8eTss/bIsZF8Za8zdN0Satd2souisxmA7ULi62m8fysXZrNB4oveG5Q+p9w6Fmsug0
zphXnxxWc+Dl/dT5JiarG0gigQexX6DjY33nmzNC/fe9rLw7+FViVBTdzJPoPBylFmokFEcEoGYM
E4f+ImD1nHIsLL/pAYKlfstcTfnGNnnf6qGMKqSbxfETPkzixZAEOEaZNJsRc03qVlLtg8DX2g4e
Ju7XNxk8Pob2R58icrrkq+uyRmDXxCLRgdyDc+eBFAMF6P9Igx5sF2JULazE0Jer4Lsb0w5HZgS6
GGG24B1u23qfHDCZnpuFUuZcAmTMOLerU7DA0on/35N3AIZjDB/ZY0Ejs81UMzvbeCWK2ycPomxP
mHZYEAi1ufx24fWlSNMFrbsgHeS5uW3KrMnzudFQu1not7aPO27pjV47iFimzjnsY1c8tQousa48
jcPQSSPOXs4vi8TiDDlRWQ9Rw+9jJRo1F/d0v1jXuxUj3hb+40b7ifK6KXksxPf/0ppQAFAX29Dr
4Ly5kufLfOIyE++s8VfluivcY4jOR2nSvmUdurSwLBq2DK3EuBrjPzeznWqX7PoMeh+LzOtTdH3p
1J8xuAcd8DY6WJCyv2qB2kUeM2b67inobWtqs3xMvzmPJwwN1AhKz36rdzgTl8TRoiongJ4uCpAi
TY6QNV6ClohDd8ScP4lHLAJrFqyQ1ypOe6VFF0OFlZ1pyMh6ldoDMWYpZj2R41niKDuw63hllskq
SYTwBIKMJSH1phZSSs42MJIIbb4BkSce/BH4TRVaqMqm6Wk23GsPhJson9NF8FRSHKrKpAE5mGyF
lx77N95B9KZYTXW0rCEZkAIHKAHhN33OWm8sdq2zdWZHYv2SuBsP1khOhsc7yjmPTBnkv7JOCR3B
jhDRAYRSggKzoAFKKcz3f6/1MPXCRjjImcJoJAEWZLFgiyHeyWFQt2LOEp27uvJbexqQVpg9mINz
buysZLlLBDuCtX8ptIOLTKoh+VtGflpspw5UAlh5uYkmoChWHLX4iIo8lyztUMVBY8rcgAzcLvRe
en1/mY9vcoMtrgiXb+nPoWBRG0VunmaXW4cYw0xix3sNDkpDAG+HbfRweSON3JDr1WCA5MbHwz9/
qxO5sCPSCAybAYSDf+RFQda+5hJmz7x4cTVKeWPt2mE29b36kkfjMadhJoXd28rTOfcjyFvD+607
oMdQXXr5v/f63b5tUuwVViWPJ4vjNfRyl0gV4Kf1vYBZnsxC18f5U3j6T67XS/ksLlHHyppHBkOr
Sx8p1L+W0EolEL4YazBdhq0T3GT1l9FMBdQBpxowKPVGQlboMWjdY69IzDkdrZ3KVGPEb653Btxd
9qcw9TXuDU/OX46KKQ2Y2nlbtK6bPSvB50jHSXEZp1KgBvBNxlK8vIVXvQTtCfgXHsjEkoLuW9yT
WdIeptFBifkc30f1fc6s930C/xvMsxPqSByrJ8XxmEGrIcczrytkKFmj3KUbgeTFSVreXJc/Ia2K
aQlu2sZQfRWzobnNp7hYSZNbunhE6C0a5rEE6r7Op0QboLHmRP90A9Coo9rmCUG8er3PqrhZOCmY
bEM0Kdvy8m5jHVkmMVdfZH2yUcA5AcWzxUpYfhw2i3F+1u4X4+qH85IHVLtmehQjXeu3kRhjCrpZ
2OCkKuWRXKdaoyKdmTyqJsDPICc+94HiBNwK3xXP87ssgPRQfygDq/NRXeQtAVynMfUaLictMCFn
1QQFDGwOy41cMdw8bgW7f/LQ9qvt26WLLiBFBabpJJBouVcwty0AHzLLyCOeyDy+VKqnqCVWxXMs
f/xpl7tvmEyNYRPxf5LxobcuHUb/Ef4IxfcGXtuEv1TsrRF6KQPtatbF/9mDHePzDLcKHvC52tJv
I9FlLBciNiwsAW8bILHKrGD2EVtA/46nLyl+bbEyW47qUJV7tPf0Dt0pQ4f8yKJjUcrSrOirQs3Y
dSL5KWBS+UuFYr2jS2cWVvIR9Xl8Di4/agdv5D0uY+Guc5NuxTGOUZXUToSkJPch+5FaIiRZI/Zz
DC4U3c4OK5Cjk0BTPvOANGb2rE973n0bw6HMzRIEdyl+wtLQTYempOBCpd025LJWHrLd/T1uf/WK
sIC3wTt785YVeUHo/UdSF8lU4zQqd9rvt7tePNI9d0qE2dgWdcs861yYQFam3+Btw8KDB9oKyY/u
Xfm6cNlqWmqupBDvqHBf/9BxR398oN/LM26RWaA7Q1mTbBybjy7lzxi8lPlfpCTsyPvPtoKhwlri
3CiXTnyLm6ZcAfRsa92R5gqdpMMpexGbCkvOvOX4hjgt6AvjHctZQrtTQTzArprN6iCb3TpHTk8+
N45CPXAJmaaFZBKQNfA8oGugOP9qeGs7kqP1yqmqCWNRWd8v8jqoEE8INfS5iEKb8gcyn1t3+FIB
si8uloznOYIEx1b7tHp3C52rEO9/2Lw+fTYzm1qF4m4j/iGlWZGKR9XF96YVleTiMwEfTw7n33Cc
VJ2+nuI1zZVnaHsmUvS/xsV9i93PAw7It0xvCqujsoAXN221X+ejZYtuyOsReOrA1YnNzvjgepEb
OT4+GNx3sbCVqK4oWC2pqaCYZmyrxD/1BFjLn/n3nDw0vdMu+qnSzWzoN3ZZDAc9j93YQgbO1bIU
L/35fLi8oyM0HSYzJDL6xZwAOlOsXbHXwGPthFTcX7CySur8iXufjrBYzfYRSYjIPA53V4ueQXGc
POMsROjKypmd98f7xwtImPhx0MNEZa6J6ACh6Sx5El2sYUTz88svP3xmkpZm1ol2p4XCvzJ1dLC7
BIEjcLHiTeKY3xP7yO9GdgaGc9HVaNtOa7vswkdBTX60W7piVhzh2+zVlH8EdBSoZnC1k/ke9kd7
dPmPfJQFC39q+0NW/NvtOTAFlOepYnj3nd7pmvNOoXPk0kbQwj/96pT6e1o9TAlJrgQ+FpF1ANpB
xdw84tenpufkdfiFW9nFJ0AtF8ODXuvWNKDZJbjd7FAVYSHDOXnS6dobokXgCDOCoxKRikHHBF5a
p7b6sAbi2dIEk5sNilE8725ZbURRl4klyZN7D1CvcOUjptTswoPwBrG9ia7KKzD7ORbfbaLHgnT5
6fS9zd0Eg1z7jaDCqbRvUEYK/r7psjHE0bXNuwgT2NvAEDugyop1Qpb+6uIKVAWIZWfUrsk7u/sy
SwchkqjeViVTb2MT/B88zLQt9kYWenpTp/ONPvliYQ2m5boI0e6wtLnUPsMLdZDW4R2OebZPSJQ2
Yl+sQBogbzW8qc/Sp79v6oBI8tFCmmJOyKuWvG7n8rKs9pHzUNH8UcDca75uAN74mxJ1wwCWW1/Q
Y3xAl4hYOkI9Z7fcF4EVZ+b1R+f34lPl+daF5o4cUeFjutG9Tbo5Ehg6omtJWPSITDaqAOJaWqU4
VgNfFMnJJbjUoYvcpH59gfFjxPwB+2T6wom2xRkHNdLPewsWNBbP6YKawKdzvyKNbVzK3HFzDWWA
4p7NixqCk/zx+rhxfbqj5P9+YluI3W1S5yjs9ZB4KhLiC2K/nEQ2e4X0lkOCpJ1roNdxZKiUCBTF
eV7VFUqdOAAnlsbR/XBd0CvuPtZiQo3cn1nuRGzr6cjcdwpkKOAoFAlkbd+25rSd/5+5fIuzHmJN
ds2G04oWuRT7r1LLXF3eSxvatahai2Y9DH+6zr39cc7xAsi3l41s2Ja6rgUDjYt0Dx5+1NMdWvu5
KFduqNzgo0MGc1F7eC0B9qmp+Zbj3zgY5v+gYJdguz+BjjGMG991S2SaylNFHXKTZjRTAB55cqEV
L0KGTQYy+AmsK0AsWwLzyVTwndEw3iaEozCq/cmRqfq4X4hHfwG8Lz+5bPt3j6yOd/imdCmC7cMW
TsAK5OX597MzAyELw2qZeuPprQqs/ocEFm7RTFV+X9cUrAd9aniMHo4POW5G9SaEAJf6+5pPavHH
fJHiex0EsOCITCKsYlPmaeoC6ql6eFvKq7fPGCyU1hY/4BNsSNnSUIZ5x7t2b/xgyJou4am/lrv8
IhG9X3ANo2eLafjlTn1pH2Dg/EJudQgkrkzr1LW+aqBAhuTb8PAj5pKwvxF8H4dMfGAecU20opPx
BC5jM+PYK5HmqlJTpH5lszKlC4cFLFRnpJfw0TEh9wXe8DQo8NEC+UKlD48HFtYereYR4MicDp4l
05eh+bwLNJj/mTRLh39jxbri2kmd+Tq2d+0yzFoKGVHfczkXL1ZkGg1UPV4FmAKO+A4AMcvHMYNj
hbJpFjp4cmiAzxOxWknoeb3vI4/AAq57fhFWJtB8SaLPJEUIn3LhPyEZ3MqHyANg73jhmlE4gKfj
tF8NYSzASfdASbm6Seb2DtvB/Z7AaUscEDpX8c0R9b8moVCoz7Kf11ePHXqvdiALrreo4suqwkvy
nf0MQfH0vNk8Ss5FxOVB3MWoG/+JTUPZUXS5Gs3XLfP13sUvdHKt3SV/Gd0jzvqVoXT35DLMpUlE
aUU19rRrWhvDOEf52fnAxzBjNySdhZHADxluPY0nxu6BekhzoG+q2mYYzZUB9pd4yJosCV1t+HhG
m9iDqAwdZC3B8RTGkcAHW0avaOgZjLt+joRrSc+hlstTwNq/ovbHj3FLUvwGJnRp5zN1J9ZLMyFT
TM+hjabMOJk/4tuPDP/wSFuN2B0epgKjULAZWtkP74W+qBEoy9JoTM1TQmiGJJftEoGtKdZEAtrb
WbT3y8uGTVzreAWD2yjyTz3Urs5/ku/DzhFS91f1b5uHJjzoCYQxFItBW0oHCUZM72b9mSdff0/u
Zet6F00SAtLFpaZaRgFbcIP8PrAVFRX3GU3TzmQfP5Ermq0Zpc4EmQ197VF9nkHXPxe6p3/3kfWC
Wn1R+ezA042ojl7gcTjAI+q6T9B8+bzuPct5Y7NshYNBjjAwqBmFgDH2XqhBvVGT9pUDSjGKU6Gy
5I6mv2ZS9YddzfWKujpE1kUKWRoQiUdyCagvnzoFiZPmq91Q/xVzasz5svV7KzcYsqbd5oz9Sz1K
RfyzFa0r2CYSJdmlVNzdtNb/UpzFYQZiQOBypND0pdV7MbqqPkKfrDV/AZVji9+vSjZH4KMcNQvo
hPWvJhOuc6mYKaij+IKam/fjsC1ZEPNYNTUkz2/JLp8QmFXVUGaf8evxQ1LuLSy4W1hXKFhO9ItO
bimORGWZ4THwr58G7Ysh9VGemAehE8RXn5fdNagc7IOIWnDIT0x19VrSZSdYfUWmlNobEMcECrUP
r1a0F2eTSn+weKaZ4Yx4yge8sbZDzvw/zFGIk7VIGsTxYwYlEgoKBrWY7C56cD/Jm3Gc7xYMzOix
xx2d9x4WLzBqqES8bnZ4Bk6v+XxN7nQFcOd5pWst1KPnE0n3DlsJ9VJ2U9MNtYVol6IY/J8SOx7t
HPuwfi8g2AmPYSyoduqZ5H1buFdst3iGORLWgzUPFbAAzFIwA2VWb9iV4xEV3NzLUbRvSHiigFvG
lQxEDEXvHQcuyQLCBVNx+56KqnGMo28RbMiN4UpqEQo2j1+Eqjl3QXimRqfAWbjUorlle81wW5Tz
OfJhGoZhsNH+iN7TddjE/nueRFmbi/BquJMGj9sP3X83xmTPHenXwi8rtXDyh2vILyPGsMjR+Ifl
Zw/S0ctUTWIUP3QjrCHJDDe8eqPVSOzb2HRa42wD9ysqwpPPn5hJB7+sdkoLqPAM775PQyqoxq8g
A6DWmJ817FYg4wtUZl1s1RJBsB7RKq7sLTfAE777EYMwd3ubrXDrOzSlQ1jFysqWs18un5z17H49
DaaWmWH1PMQSFaDQ2s1a1DWJPOVZU/x2EjV5U8nkWIrC31dW8gx2ggbhri9S5IC+C/l+pOkaEcmk
jtQMgaoGjlGxU7LSASInmJbXi0bNd1BBULA0gr1kTYW53p2z0fL1i6Mg/PdFmT0rENo5skKEVL19
y64xdC3yMQ1qe0FExlDnZlIuMkKqK5gKhk4rupVKCrjD83ANeOVMr7IpKyGevLsaHheZDMVcIKmg
phXe2OU1lRN2i22N2YYgi3xdLs0A0JdsQVGVlJJqfr2DfUmM01Uy1yzrIszjnJrfiiv8DxdomKzB
cUrqVkKSLBsoDxxLZLyrASQw3FB0KgaIml8QxsEKFj0MeZiqOotllTFnRO2u2tGHiTGCVhw2Gde2
pzGdztY6oY2sA9t4ShYSh7i9Bgjv47xPaPFDArqNSjXY+m0kugWGLu6EI3iWn8xmmJdvRBYk5CaU
wcnNjx5QMXDReCRGOO2gjtP1SseK/nGc7tZOU5+FCXtkLe9M3T7WxYtRON4BRg48ImvqePz7JLvU
O5lYb3R9t1F8OI8JIPjGxSqfkqV7RTeNhDYNNkvVTInU/CWwMFu3wgd1mbmUb5vI94kHDqq8j08t
bG7wL9C0uEQxPcjTshWVv084yfoviXQBp3wuohy95vRmIr6nvtduDtfNQ5KnqA70lx3ypX78WQES
AKD75lYvXbIf9mSXmjSsxJ1Cd8Tdu4vFO/PWJvQVNt+A3V4kAIMKzlmZlIlPQwjxu8TaSK5f1DC2
RdZzo9L61u+RCfzdMiK/G2gQl3hvb+grttVEySjHQz2SAebisjWbmzW1Xl2pLmwTZE7RLkODrOxx
BSmulJvaeQhmBsem/9St9PwKVY7dmh4K1+SKZ51o9QUcn1L7/NNMRHeD/n3a13geK07x/MhPrO5h
kXAxBS0aULNfN1+aSZalQpS0OxPU4Ca/U2+vWi0+Y97iGHbVBih7MxjggG8JtQ/M0zcVrPB9uvJk
gmFfsoORo5WDeyr+RNcXETPtiEEknKl757UpIiK5llOwtMFpAxhrr9Tn3j4eEtj+8cJxxntKgrWF
EoIQXZxDZpNetcRq/2UBDBbeS+m77QKtDzT1oxe99aUoIo0dX460Ccn8dTFbbSlatyxPb1GWOV63
nbNwcrLvFVaNslhSvyWlP2/cv7D8hgF8KujVCMaBhOCrtwwDFXAASKw/CHfiKUqUUu7ZxjwbSDA1
YxI3MQHHtlsNrkLeRUPb/sMXSQfc1fuMBPMOLaMKiMgUSW4fRXxvkHEmFM24CNZVLmBl5/9LC4rk
wp4/3zGloqrfD/9p+huRVrRV6ENq2zF8AZDhqDhBGWTmxU8XNRbe6dG3i+z5BnWbrshw3JCmjf+F
6hAqlwBJ/eqrPpnKcbDn6wq6cO1iT++S+w2nPQlXKB94RBlIxHc7W+Rq7AZP+fYH14RUy4fX9Vfj
O/hn6e/BDVtQmFoQix0gSoFxntzovU6I6H36D1CViNjq308Ff7MFhNkufmwLaXg/BNkuOlWPTZK+
oWg7hsghNcVd/bR7QVdXJmH3lYykmkzTx5gjiH5Q/Je0pMIh3xUiv8W4MfppqEAm+FstXeMlwzAz
yjZEpFG/9tqg7Z/dgd7pZJQu8v3ctVER0qAj5xMXh1mfbFwVJLxu520Uu6Eo5fT3dA6mgrh49jQl
D8L9Xr6HYCu3na5roNhpAGuOuZboQmCL+afhwJyNdYP/W+hFmD1AVQxraSjllYnX9gYMayANIHUV
+2YVfOg/8RaYKvXk5jao5luvuW7lBtc9yd/hyRM+n8vu67LGFQl63oQk3weQwJZQjnVOcg72JX/p
P7D62mrEGWhUB0EefqTesc0xKeyWjbI4JfhrW67IViOEonZ3rfGF9hMdC6b0Cv7lL2LyC45EGbxp
9hrN4qp4tPH0LL1koxl0ncOnmhsa5FwT/M/w6cs6/twMvJP3qPXj4MNhA4gBBOmtXFbZAHW/iOPt
wqhTU5SZhZ77t3MrQEXMvXDNK/ySS9Ii2HfcyoI0PtIz5Zf4E+LsZtr6UUKy/tzYF41EZ3RLHoo2
bFDwKCQLSWuRzKdMUHOeepZ1W+0ionyTkbQS5FkWCt+3FOJaXa+IgeFQwDggOuOb4LUhtDfCnfid
10ceZ/iCBQnE7pCr90SwamjFvzorwhYEdRwRoEQH8Fy51OAnskEv8tnF3FPtQbH7yXEEV/J8+2QO
Re+Yy1Xkyt+9NPu3Tv8vd8wUHL9Re6tHCO0CRbXvRKmOgRT8Ks7IgFQhrCL7mmo45NsqoEM1K++1
7PqDxu/CGpSSWTUn0fLjWy/5BWp+NjyvR8KVqTlTQszgQmNUvX5EJvG4WJgAIG/SdvsLTNUgm7t3
mHC4DXR7ojzSjSBr4jztT/IFK4kfD/J7mV+3ByuNC11BWhMfrMwZ/5QH6ON3YoPbFh8xj2Mu4F2x
Jt5ZaIahH1SQPkt7FY+uT1C6s4WO482BXxzrFZi0eF0KGYnG/ch609EoMvVizDyoUAVVMUYntgpM
JFi9DeRhyFieul6eOu/t5532Nhuw6bWn44O+XbymNIECavuSC6UWZsbldZOhpttlLM+vfpC4FPTi
mdXSD/zpCB9oKpyrTYvrL0vEWEBTMKfBRYgl6+sCFUvqaEwHaSBLv13j06ZZCp9W2yQ0t7DwDkmD
CkUm/76zwgF2PXV4KbAhfImiirJqwBrFu8F5c2GbnWc92BPLMTKrRMcBjDUJWiMZ8ea+BtziMp8s
x/vD4pvXfCD0O2NUN3qcX0st8SaYrB7WLnHSW67sAUNJnH2DCjSEPJhorHov1hJ5xL+k27UdAJR7
b7L3obnbHQ+wLp2TePL3hdc5e1GHXu5f0dkOMKl9JRKGv9g7VQcDy9MrM0A3PvjhE2F3T7/feSeP
MUy386bqTuKH4FMBmU06exETF6RR06Q7v1+O60vYqnk1JMSI/rgnYRkxULeiSOT0CbbtVuuUWYIE
5x6o5n/oUe0HCLBDiOioXTq3hrtNuO5pJqu9bEIqu3+q0wvhktVCOF9vMm9weEXjd/4gg7JIrRQc
c0+utaFwBt1eV4rQkcDlWA/RoXjM6dxE/4vj2YOpjK6krLcGNVO2dGIzUQ48rLOpRQuJ1tYfeXYf
fme4KQ9d6x4Vo5+A1Z6j6cRZnWI19t1NjFxU7s4bHI7WhMO/DaALOwS1OF6qg59Yl/x9mAZ6OxKB
yXpG+GJQVXBKFk6v/vxCxHW3W0K23ifN4FBDfOC445GXFZZDeuFEy8NF0+TMOrDvVlusN7sZNEcw
6alyBmBSb/tbslDZ//4imifv9nZwiS/fnQgTBB720eh2SZDm0p1apLjtjozl7fWMCDq1qjStz2fN
Na+cIjL32LUwBAYUj7K6Hma9vdCuiZK//5IxmGZiu1qH+9LrhwITd+ukBA2pXZTIu6bGAeQ79MQl
WBBVvI4Tq0xlzT/mbS0LbA06uGA818fFKqOdaQfoB5fXSneBn5+gMr3J7EFUeEhmEAqFzmXtN2Pb
ZdT3AT7Sfm/z4WFWlIS2opuLLWCMGpSCiSv5isoDcyB52F7SM5/ZmaVEnxZxKIV8nvwsk5hVyCbC
QJS6xSCeie8nBXIA+aRhF6akqUmrwTBukVASNnqHwyL7AZz3RKB0jIY4hmhTJ+78w6zS4PpXvm17
ag0ogDTJSmVzZqeIKEr+n8bgrqfsRNtbqSBjLi7MRkguD+7t1Wuii/9YQYWRF6iQd2nOA1tfy0ns
pUjThflPUYhGb+Tpp8ZwKLuDsnYffxkjawt31psk7mybg5ILF++45wN+611V/XErmHmIT8ocxlsx
UX7MWS3gTEnoFpccjsK9nt90IAHMWc+AXWw9rjXSr2EAOReTBtTWGZ++2e4wxYARlIktiuR9UA06
2Si2JbMR5XtQzL7RaK6O28iz/13wCpout+gJ0vw5WN+Gy8cCcDz25MkV+bCA1Jr0xEZp1hd78IIV
Xdg2APPocseTnrS8kznYZKQsAiWsW6enkSWp7EPRnzN8BLDwl0u8KB+QH9yjCO2n2774Fvs6o1bt
WtBCAeesjotafVws9mtBe8/oZPITE8aldwS1UuafiLL9U8/NQ+s1KLiJFRhl3z+QBzNa3Uxo31YE
CQ9xuIT8FXgaO5ERikLBJeh7BvIAewDeFaz+zj9Jwl3Hso3N0uX4jTajqJOEJWjFlVPPSszPc4mZ
Qd7BKerFfyqHwQ87deIyhmtey2bm63EXqgdnNOBocGwvxSW8Y8blxLynD5r05ZBaGyR84Ax/x0q5
9Yw/0stc21CfrZAxWGcmTmTGpiaVY/u98K9FX4e2RflDWATn6PzapaKXggWB/XN6v0YeP0y6E6ro
tEYFFPV395hVyGSBwIMgqMfg5qOyk9tSrgIRRBuuXw+uNq24GHbSr++zdFiH17RzuKVbnAOBRu0+
QLxX3GHtoQeCUxawX1aHIkTpmZBygTDUvU+nbAyyIWQbnR3BD6vjFmUn3Xri4DO+uWWN+rwesJGy
YlkJ3S01DQDWjaTh263AbH51ySBJ2JU1QrsOYV/sUBphm75ybK7MXp12GlI3bB2i8kTIqSN5+rA8
S4NqgdI+sVDSkPk4vxQTHn8ReSi7P8tB7FC3Akr/rP5rRWmtEtgflKiDLy62sC0VgArJDDeskz9W
NkNEJepVwGPzdIdzznZnoONEjHxm8Jd/X5WGrpC6jtu+71Vs7cUjjioZHA7vgb86HDu+rpM+WY2C
Av0/JyhajW1S6sMf3eWbN8Cyim541O4bEQ8mIEoVatcoDQPOE+AvY2wqdQZ4C0oJWYJV/iDGG+vn
DTeLNgBJvW2pOe/20jG0BtvIohsRqp/8PL0QiEh1cU8dJXek99Gdna7PX7pVWwE8lX1lcBwN+4fU
v7ksckDaM2XOzE+Q3NFGKvY9dHbzRaL/mcGmkz+Uc0OeszX/vkLVACjWhcXq3/pLaCjD4TrMZUb8
93Hx/8k/PuxMIYYBHzX65K+YOrUxc1xmOlbuB6fDGWSBWr57/2k76aoPCq11P0jfvtbf5/xZ0lkw
OnZi7kf/+2ZNtTTfJ8ipSv/fgB3MkY56uTFadWrbavILoyWh2r5WrXHFAVM0xUd9t4h8ccYnIu81
wzKIKr67P/RwgN3dYkSBdsNIRcCsABgtubTXHobDTXMIKnM1BgcNq+pBh0Gw14vralRrKsbRnv5i
PUV1hvhf20AWKB4nHilOs3mIXlTnYS7Ote8pyYt/TkCYsR4Qf5jUWbFpPZotSY9S2kYndhZ11oFx
vnOaL13NNoyHrMHUxbFQev5NtkMYxeUdqDnP1YmpeY94uk+0D6WfKZT1umP5zxU9sFBTgLQCu6pC
FA+hzxeFCZtNRXGAk1hXQxQ3oQsqGufdoTf+JbljL2pf4w1yHFw/Oa3wijuAHTIBud7b5K77z8J6
F5T5J9v77bUEVkfo1DJiscs26OgiD9hFiKA9oRldXDUdGFUL6aV1ZN8sMxHVCQBjbZEMRP6FPUZN
Ti04xK09lqGaQwQKnHSNXim+uT9cKqjFdLWOA7Ha+kj1T35KT6ne7uAQAoCGDHN3Mbny9SvtSEx/
i4uCCPcDT13OXihEUq1NIzKq0HQ3xteyAk9r/pkPrxH7DU4jROS3hG2eDLQ4EYCzTIlRPXIUd6QZ
Cc5x+aRfYr/KDhGxHA/SydVo8GB2C+BxQnKOHdPK1/AXRlx5Fx6VA7wyrL8DOCATG1nKlyljVzK8
PDtc2qvfPqt9KYKNbN8KFb3TONWATRFZGHY9MyouPmDajd+GsR5SCyDJMO+SIaOxKKQbXUo4TF5M
dUsV/OntWdQNPPYsg3o0vLAsg0U6JXpS+awyZoe/eoDDs9+eM6ya/+LfVob5zPOIVLLDl8/b6uVm
PUBs7DC4zqOa+BM1pmncMzhBinrsQXcAnJtzEUCaVWtYKxwJTQyNhpPmbWvef+fiT/otQTza/jvW
fQ6mSegnhjKkQ5Str/nvqUqmjEg/w46B1VUL6/A5siehpfYLxMnFTk5crpEnM6PpEWwRnqkvhXB4
YW66Du3fgOGQpBtjjLLxazsPyjkRuNSFMFvwDrQt5Fi34MsqoqijDrOVs3U2daktxtKvs9/XnhR5
fHyvqhUdKgSV6sudKK1pXTVnhYVJ2cQ/TbqImpxVTZouPt9KIJw1pLKf4ClUL0JG6PyjK/4MvTdy
Rbyc9Co6dnvOesDLAPPNcDUaX+X82h9WCr02ESovm3vcPY1lbfyXxKJ3IQe121YNWiuuykkASFl8
wsx3V1Ry1e4V6+3kCox8hE2Ql9iAd9xUDkC8zlz1k919uwkZFAcj4/tnVpqwUdoZc1ZziLXoTPDr
Z900tYgSDSg2OjxLRwLNGz9X0B5H7ROYxK4+fNMvZPhcgdr3PsiFlyeNSmdiuaYJYRbemerE5vTe
zq4r+N2WXn/Aty68iJ1XUiFPITLEZEMJ/5OVtuGFsugy87SaXK0bP1OuAsHtU3nPTtz0vRsweiiz
i2rLPikc6PP7fJKOI3dg0X/Rs4RMJfuh8Nz6Xii4BpOpf7/5j+Oz12gFagyHtzqsoObFt+zQRW1J
ma/dz5US9CXBrjgdQue5D+FZobnCxlOZVajvJ0dC7g5NcSNlSQED9vwSlsCHFE5gYkQsI30APjtS
5EVH0q4kSGhCDi+PE/qXc8kKDvQO2WArN2eJuOfnYGHXNhbyQmXHAe/Vl5eOHJZlJ2jai7zsnaNw
wn44IW07jMWiwUFkfG4JeGFB/vpPm4SxxlbrYu2VoztWEO49w3M/eGVkFZt1Eeqan8ML9dFHuXtT
gj4mOoHWdAgWukXel+/Z48sABIhs4H0YHtbGrWXxM6NDMx4R4mTpooMWa+APrdPJ7YByadRKL0hr
Gw79yaKxoCr2q+V7IME3i+gsS4BCAGZ7qJeUwLcRurDYpxUoEFkUpjEHfaRvMTGnOyT11azj2jQy
v1b1qYbjgtx7XdaenTcVCQk5+mTqOpywJhWPXJ3R84ZdHwOussW1oHOPRpklAgKyhk+VCyxPqDp0
QjSDYey+rYBDFLfCqAQYk6fYzWz30C8wBK7ivus4uWxiSAdnJmqRWyYkTf4YRCb6lUSe9rWYBg1M
aJrKz/B61PNFSL9r9buXaIxv6Ho1MglErSYhWEsFzLtF/k3iol+xvyk5dBbmYKIs5mdJ1XlM/HHg
wJiINYeev3iiayC9QZhfDJQZz2qWdVX197vCB0FVy69/kGQj9HwuPkYPpdKkdluhfEVpPePBULZ0
GlNDOPBNdzWFM/kb+CFReTzTZU71mHJCkR+8McmpbVcmfox3NBS4qphJQQWXVdQVCxRsi6/q4xL6
ZPlqjy0zSxJVs+BuipQQfNyLfHTJWkY2Hj+ZfgYbVLPvkPU5wATjaxokwxJz4zIbImu9P9kEMjsA
ne69C7o4+kc871BMav4lY0b8foqBe17NFns9UZ7lAtwZwWYSbVaP7KRw8RbS0PNDzq5uwCoZMBEI
x/kuKCWDyiJ73JukTW7Z5dxCIYeNv4ZwNRJ3p5AaoPyjkRdD91em44ahHFuKHOtF0P6//TqsEZGh
B0YItU2/b1MFsOegye+B1zfMNnXN3MtrS+sjPUgXSxWhlObl/zwNTeDJpJdTlNJNsJx9H5wIwSoA
LVT9loSo9ZepouwL1m+bNEGY7NDhnomxjgUs7mPhEmV+DcCpdRiaIv+kalRSP3dzq1zHqmjBU6cx
n+LzNkaRHRoLmSut8FZh8BlF7w+rvHW8OebKzTshluKL9VZztNG3LB4SF6pBqkKE0EwaToK4aEgB
9xCU2aSD6BCRyByQbTBZhyhKx7/cxKgnx24LHds4U2J4H1Ajw7JAs9k3kZg84lM+ZfQe9NK/KY9c
l/3Lrnfw8WqhIaumUXQhM5nygFZCoTABbAl7QAF7syZAw4Uadtsymmsolw2DWcy8vbRCE+TrZDUS
ycHufW/BN028dhMP/X8NQ4ZG7TdAWmOFGTHM8ibIVvdvpKv+kFYlOIP5qCt2R7DuuS7iMUIB0niO
Fzfier6jhpgP75bgT37hezrbhTWe00DPzj8/vffEL7N9CwhuPJ+NEiDlvBK0rkFhPOVKVPrykD/t
IOq0bWJOpbvYwOflfuPRln7TAbekKr1j/jnlzfGoEVF7F5TpI26gYzGvmD5HY4gbnZxtory/CxKU
9t3UMJQVM9mkyqlAQjT41ZXZkv5g1E/uB7EAW5Oc4ybLFl4OI4VfLqMffCmORLYkqJcF868KBZKY
3aprTQpsqiBkitCVVjDETa4gYb8cEqlqCzxJfdNCsCkmHTcolw3phwhd4/FAJQG0zfwPm3HxZOmD
zHahx6CQmH2EKuWtEdhE0qRHLibnqJ8xd9ifSFz75dQnntaEdj8sc/JhKrf6+Pq4uU/peXng/Jl2
5s5cwGrsC63iMLLJ73d5i92htpzSEY7YFv39K3DQsLMFXnwI68ZiRtMsen0Bm0j4HItB6T1BzKzr
9zTTuSnAUzY3TlvvpmcmFuZ8cNxCjgQBIzJsLQZ8LSgGjm1F3LVsMdVcWio6lSJzIQ7enr/n4Wl3
Lvu6W5aD2pRl2ZtZztdBPFl6SIJ7F2iBKVcav9XEW1pOYOyK6QUmDmBgw/DV+Fe8PmTZmB3US6/K
+uqvqQ067O1iXwpACe6QEwAsiJL6bivpEO6yRIBjvmCopaNzAtB+YE/C0RHhtIwq1H6zfqJqz7vj
lrtJvwkc4ffw9Vcc/E+ARTW0XF+/st7yLt3BWTyaEUo8LUQaBE//LXEZiuwDM9VlbW3EC4ukfd0V
cotD1FMluNdiFv19/VKw7craA5GPicTXw/edJSNk0/tLQhgzJFhT81QaqvZ0/SZcSk70BfTOpmnT
G+bsERm3u8Ub6OHMUDPf9Xkom3KNUhhoZmRzJ066FqmGotBbjgVPM5SkaqzS1MIkSg25VUm/9MbT
BN8KzlrnRCuKsyndiXi+izFl0rIOI0FgM7VBBzEs5PlupXsLFTW/ksU70yDMu9PLaRGTS7BLrjzt
3i9M7DyUqjYNUIxQU3nmIhb/OJeth9/4UVhLbwDwJayio4vpEW2KZBLdeuU3wFtLc/CWPEvSL+vd
UECfNiT45zO9ReoBegDWOYmokF/K9usq/NU4aAPGMZBIorjWiL/mFE1hW5B6l4dfy/35HB2DszEx
+pkZwUyUZqwH2uL/K9pLyuNglVzqr/GAlzu5MP8OigUqy+KgaV8Ubyb9wztu61hOJRct+Ob6OdmT
wEc8/HL+OYDYI80Sll2Pr6r/G2ypvpL+ZWq2dUEMCP+9b5pJX7XukmY8zoSNe+XcGR22qixVhHcU
LoJnVHI1uYu2L+ZnhxEgox2fz1AZuNMFJrpM5EawaRWDfXlZ9W9LTn5dGWoCzzJ1JvsGsNecSfk3
o12p/eUITkt+6sUU6s38U6/fHDUAKskAko3EBJU42RRJhnoLzASCy4TUkleBag+Q1MUBzr5VmXM9
pbuzk2uU96sC6bwPC6yt2ER5yG2uY81ExpJ21TawGHOOtTKbFJXWCAZp70k6MovviHEurxNxmWE7
YAGPWwE9x1jCMJ0GmbWOCvxpYQyB/BGhCRi8PWUR4I7gks6Blp6IeWoXrHrvpqINQf919tLwyieE
9HznieES3iHzue8X3mhzBfvdlwfn4f+jbFkuZ1GPgOiyO2QT8vugv8btN7J6cEuSbDbF/ifYJCTd
HiXMbvl5iqjU1MjjPSfOmnxORg0tkfW+wVPiHbAsi2olyU3Dv0igOdNmTqO/eaY6BzIRa0mKKm5j
WNIxY/5q4sGY5c+ZRLuSOZs4VXuhlYGPzmwKyEoz8kuiJ9nQNnWS5NKrrHVHr9uYrhzX2Z/lK2WE
GOHCYOYY3A4NpHtYd77WxFKqVZu5a89t7rF7nZCry+ZYWAg57Lk7S/r2aX6bDNo6slvWJMz+tluF
pqsL0hu9Ob3D4uxbusC7qTr6uC+RIsfMavQfVrJ4EKbbBiLngzshUaTgaXbSg60Un1SneC+9c+Hd
oiODn5RA3R+4iyHegfPedxgP7vkCl4IyyCbo1lD/fPrdxKuWl345vrGzXz+rJMI5+d0pWUCCAnvC
tgPZIQx9uQFBmd1iFLpn2eUOJkt+YzwdOU948i0d+gZ2RAAgyVc8KVOnzU66vAi7CWJZYfdVKoZw
uF5RYh65IM+65VfLXGutqvP+T5uCaQ2apGlOQA5S+Jj89S6cp1iCdiUxL+61h7Hq+8mjsJ+rHj2c
a+i0CFkEVBy6BVqhVPVQ2yHfqCd96BbXL4RYQpCNtlHvLsXRsFll8vF7fO2ddGcrjIjZpjDOPKHf
xjv9kPhTGyeVUgDWcWa0mW0v07zoeYxk29/E5dRFHJV2Ejv/Hw/RUZ4VWohF/wreWvA6r2Gw/h30
gg0U2GSP3I1gjTg7ZNwUpyaIlXUvwI/D9N2b34jv6bsrgPAlhw2qxnJ69nRnILJNYfMEL+iX44BV
JmfKVoViiJoxTMIT2Zlm0nCEU1tKm4Z5Jv91aYSq6R5/mt1aJfIHGo0L+kDdSSwnF8YsMGGFJQDJ
gwy45y+/zN9Wa4GohXwbHggJuH8ubXll6xH11hAgqDcFHzcRC3vVoauvL7Zq9dfY7xBbdA4Bab/8
8tg50RTi/QyI765op5v+AH8w+fWq0rWGnIUwN9c5MSlCqKekWvsCQyycLXBhu9F0+pB8TY1tPQX9
10SbgHuc6oh64B5RiAz8bIbk5JX12yJV1PcbFJdl3QNFDOFHFbY10klaCOyCelt2J9RC7wN7gK/s
FqM4QV5gMk1htXPtF5y/aHv/rt3VcVEYdFhzTe2y/Gor5/kwonQlL+6cS9NNUVLziMTKa2fjVdba
MFPpnL7P5SO5MwgBzAwbD2GM61PfAzSp0C29lo36pAADLj0b9scCL9+tyn1hcvSOuOQRImFL1vci
4PFcjgOOinqjXGcned4IN1Iz9AAH8pJtxJNNznyNm6IUrKQl8z8SAFIDpGD9dnBltx4IqPtLUOZ4
jl7aDeWf0ASZdH3bnqvVrIkUxpRZBFP65ZN0IINlgpsZvtXuAIoA+L2h2Bv3nGCDcoe/9eFRQsmg
SX2D+A210FcY3KBeUnh2XL6woUeVZYN7IpKhba+7ygzfjxT0oPtcddsd6+iDct+25CP7OLiHgXe3
Rq8NJntCnZOQh3zYJZtwKw0581DVtX9/kx69Mruq2eETclpPsvZ3HKlAXY8gY2SchslKgiQ7NwXl
clOEkL1MeXfgeP5FOtb4nAI+2b6SC1atgJR2KG6DEJH+3Voj2yLcTk8VMG8XGw2LGiTU42rB5YNr
aWGB168HVdFLerf8Jg0Ysgdo23DJjQHNN/TiehU1l+oylPNpQadeJZGXhmSFC0atsIcv/rSFKjhb
gh3g2mZWUm4Mzyl+WOxUYtIYlE3IhVkpT1j6K4A0g9+S6PJx+29MryX5MZmufERl6JNccAX61vDJ
8DOcBB1VYkxS3FglrendKKYMAlRxV4rSBWT1qRh4W9ifAix2T7EHceKaDb28VjZb83R5WUtNp7GQ
nSgDAvHM47kFDzs6QGls3R4Vrm7w1TZPhy6tzNXPFL89IEwY9KEPnm6vKtlMnjhbp6FhYbQC3gnK
I9AKSSy2YHCGjoR1iTNj54XeeOSrDUZdqUQ6cd8kzRTMWT0xLlcI9aULjDoPa05Xii9dkBVwAHHw
eFR3byfJVDArhtiVijYHvlfWdlX4EKdF4NMYMww2yBx+Ue1+vRg2oohAiVb1QTSXE+zx25ANHWjj
L/D3AnWdPmdu+lkFUAxiqexdIZdd4PWYTLay/w+KG6Aay2yugww4gQKzxDDJtIAvOvGrh4oGIN3Q
JIl0thc6wx/qOzPzp+D+dTujbKY358a+6WC0/FXzmJhYczTMW1J2YX0LDNSFp0/zubAeQWD9MBWU
9v4KeSOqDp4r2++IVcDPqSWPFpsvfJ8t6K4/tA8g04UVrSeITr5qF7wBuS42tteL1vHTs3No/UbC
25Enj3JyhYut4/ng3iQ+f76JP9Gfh0ZX7CZlwzuZjJGKlWtaHz17VV9l1Ov8PIZMXwCe2EKZ/uAT
Gnti+3TZ6SKtVb1uKgQg5bqYRJPXMritrGMAfc1PtgXuUFYTWU6D7mHX5UncndWVFFL1RWKEUJeJ
v4LL8U4PHG72deKqoLyCwpMlLzD0q0OlH3MaPaSiMwVdV/OVauuEymUMrlJbJzaF5iqALyr3XwlL
PgY2alnQne/+77uFcu7zECGVvZkgHVzmIDkVR+E82vboXgCqrTsnO11IEOMv6KiucNIeLTVFxyp9
/xJzSC4pye+CETPd3IxPNARSWfFfJVipIUQHlVyirtvWkBZMxHnLf+kfzUvX3dempPqknmUiWMzv
7NhCsXQLqUjS4192g6ZC6mixUumS4ZCk1XwSS3CDpn3zOva9hb7ns4wbaOUiX0W6NXwoIc5gK4SE
FiOV70/hza0dV30W6VZlqRBHWm0FENKr0orLuIYGhAJHz1PhufRKU8rv3EkCv6oYBxsLVwuevQfj
pFJqF1avGlHuibo4nS5iR7luYEqEc6VymQzrht2ZSnmMHoR3VQ24E7uquocEY/ZLbCunvJCi9LYb
DqAN7qVE2PIc6UWoJBs4UlKT0Sh2jNp/Z917Urbj7vClNcR1F68vdxwkUcOQIDolflc0XBHDXHc3
0a4gm4Nbik3uyXUQZrjWLnBXq9Vi/4XPYssxCsiK6XY/vV5Qy6mcCZxIuCYCwlwCAju/cRcu9utQ
c3wirE8zmrUvGaSEWpJLMEwslNLZpI6ctA0otqVotAG4JtxOfPTFTd/gxCmtafA/1oCHH/z0i+Br
bYCi7P+MKHKW/9lIV7jXAJN0J5WDoPAUnnNQpO9NPtqC6sp5WMM70ATNp0V7RgNk6itfoOx7WtEB
sLhT1QBTNSeJfp+/uDeewsaGTRJZlG1PJB8DqYuUrTx+joscDdgDQsn9YWbs82Fn90DhgJhc7d0m
tjV0YLJt/syxz7wR/T21eUprkbYAWtqP/UbeZ+190HcS603Olt0TPmUvGb97qhRate6iSUoxy3rv
l8IY3rabAvcq45H8iQL6/XZmNApLXyhSoEYHxFdse73jNQXGEZ/DSM/SbiMTX+WyBIvZXcPUVp2I
+39mo8BoWBWZtv+QAt4WqGs0al/XJU5RZMVfB/ftHSP2HuGtrQ41Aaaa/ytCo7nFEJLlJhLhAaSk
JSRQHdSQWyC9sHz5iguOzPeTYl/uKAW5IkHrvbs6vRYNA1T4z/3J9MTcgwewh2v6mY7RTqsi+NgR
NMsITbRjSRRaVA4G4/wbd+F+xs65otQl4TUf9e+HNTTiZ6OdWCmX5lbGMOLVvj69PoQ4aWYxPJZb
thlTBdxDE1JmOs63tL4z2/INJNDFbHq2sGBKrNY6B8I0M3NBTvjIiOu4W+A/UNAPg4XoV8H9mhOV
4kU3RcxPCR0cNXWNp51tp5s0ICVAX7SsKkOvejyhb5I79VQAbGvv6HUEabosVemh9nNNbJpascf5
VDdvvGvsM2Vg+wnLqIBSn+oBhEX572MRjkJvnKtqbRhe+Z56TF375UfUE1QvC1kHDpDjRLzkDav5
CkOgMPAJreWehki9NbYmqNTt9GwYEOALOt2vTVGKmi2Z4i9emUTJeDRiyh9l6Wr8iT6iGaIV1c94
Wdo9RAbPmBL2JyT0Fi9tvNFG+YUtwpbIKIY75+azlYnG/G0n79VOrZh464ckbXuZygSK229tjroc
JHelrd8Ms2UHef6JGvPFw03umngJCSoPDFM1J4obwEgwfF/acyC8fb3WpQzZmYAoYfFU9Sv8cIUU
+WhvwJnMaDZ0pHuFY1M/nRMVdqGmdMhHU4+98pXd/sjg8QsPKHf9FK7WvDlhy9skjWNbrUiqRsjT
9HHtdQolbogOvw3jc33SIuAkwMysCBfWicadvLP4Of1oJ2fRfN1msXm5dX54oX7Rf+6PTBLPoFhT
U8Vv2cDpnsE8bUDtdJ7vwkFN3I/yKYkECPSCXLo0a1CDK6XmDZdyhiI0ITDFQMlxeKjekJCCoDfM
qGV352igWy24t18Eo8a1LH35g5hscyqQ5tWMKijCE/5S9TgiVEB/OZ/5uUYfbqxyXHT41O1sT+J+
TZMdNV3IELWyEZkGn8OldYIQL5TjR3DMYXS/yNv9CuORipw7rjwCVv75g+8u8rkWbsf3/VSutLvP
BRIVzPGU04LqAZpQBI91IRNIAQEjeumARGnlBoaFbvmwmeraiKmMnmfqfsSR2eBOB2dcdrOX4zUT
zDaHKcTlAzlCfTzS2zXIiW/LqZsDIWl4eyNT5TdWBbv9UihKu9+n5R/BqeLIsGVvDU6owa+0kkET
qE3JlsZa1wYvwuB15S1xteW+Pak/D6WvxOe9svFCQMnwup6PMNhgt/v5o76kl5JMLbNGzQFHtlcy
MR5K95aWgo3k9izRakEJHtk8fF/gytImVKnOfiD+J8v9f+8HTI5eMxH0WGHuTFY9bEqJfdrlMZgS
pj+mYRe+/Lr6EZIbCxTtshQNQobwO4UohBU9f6AIeTL6808Vo9JRGuNdxNyaP6fjyakLk80VwD82
SkDFOekobxM5Wo9wrJP+JwZBDvkzBwlcqDfQ5Hhx7dU0bOAe1fMC20zhDQvqotU201N1lMt999Je
1VIX5Is1aMQiSLervTY7pbDYHm/r2XqNR8QCLTOP0OyDpcHDJ4TX12nqMGA4tLm/zXDvbpWHyWUo
YVgHczADepuaCfhBdxOGI2/msCP631YDcucDYQ34iAvsZEVYSkVCyEUZyw5BAj9qKA8PnmBWutig
FQeAPyOJIWCFuYVD9mo3DZGea8jrTygiVCysJAzJe692tmUUf4EXalCfwOeivjC/cy1zvATEHCUC
VVjrSkOoSDSlJzonEzA/Kfhy+Mzkg7W2GUOdgiOCLQVxcnrabzvkYbgTu60Jucij7sFEADTWNcG7
7Cqgsmz9Bo6y9j0BQ/ebmyA8niYL1kjCz1KK86rCfjadlIwJZG9+ZRSSFvL8FIO+Uy0T0Uf+LQH1
U+iDpNxp4j905RfN9NjBZYEyfWvPfSysG7ukfqNMlOIzb9rgL5E5A3UrWEEjvDPzqMKAlIqI2k1w
XDhN70mhNd1f7tZ/OJWganaAPaO6bR/Uq8F2XRZ/P5A5OvZOkA4gEjzXVO5piwMKj8FA9WOFwC6+
m2qlPnHUVGnGtstU2wrPOMPf/fkKz7gZlkD403cLojhl/Nuwr/EidnrUoAWL1siHJDaxcW0p4fhy
5vIZg+VYNajKaGMtqoNbHAV5QkqtXtwW+sWdt2GFA3WKjYmKJUEojQ5lOFPiTdkShJiPWyEAWyFi
MqlMMieAHm5hMEzhMcus8+ZDikfDb0Tg55/oil0Eo45Uxi1PuJEDAQp00OGUNbHEYrjAnRLAQWPR
zIAebzwE6ye0zk+hXIMgMYCDaK9TcwouftZ+FOJ1GTfZn3UKLuUpCkxNPlUQOif/C9o2dbYMF8by
BIQB5WyJG6Gdhe7njN9PROQbOX8D/Fm40Duu4wty5DrlA1t+AXIQphNCxYZE2AIBIFWMl9BjcSLI
AwykdzwxnUopUETvWZGnBIGigVHSHg0e2P4J1sMxv4twf04yXeAGRv6FlBexQRB0ZNKkqiruV1AC
ien/cSQMaVnSQ4YdwVOu2mjVq9O4iiefkX8Pw1kADRo+V5kjxkpHTNwyRtgLyqtY9okGyjmPAYs2
M8uk4afoyJukJ3Njb+yyI/rxi69S2NnSDhToNeWX4DqqU5MzpaFC+Swsq1gaPOd/RWD3oRLBTTAn
yVVCWm/kKAyDs0y50wPOaZowg4GXAirIUq+YaCQcy+Co8ACQ881BLv9A5Zh5Dxtqse4pafT9nPA0
zNUsxDwgEexDzRcyqjjlw8JhqbO2bCPRRJG+pHcYM93h/c7BeRhQC56DRrdMfnIbnbg5hVC6cY8A
3a2HSrAqzADb1YYe6biSNseIf/FprQiZYlFbyplMH9QHdVhY+NV1ILq7yT+LLeR+zkFtC05DWKtF
C+QvJZgnXEGIWPB8uSQubZ9HHDvpp7mvupG/AGMtH9QyG5ROndFppvZaJM58aSEjURc0InyI+dm7
4bW+d/eQG0nFoBQZCzCO49shK9W8FxdutiwQZBriFOucOxna5NvARWd3ZtvQW2jh4Fc/MVNCJQRx
NQzH4tAt1wTstwQAMO9dd0NATKcNdBESCMQOCcobtoGFIl3l8xPVQ95tpJ48MIS41wazvPD5Xvea
qyIUjLtaTmx+VGuo1J+7qrJ2R5Og2DxRnOiw9Ly03mK03wuFko++5HhqsKncS0tdHgXPrJbG8l6t
b3l81rLqPjGY2jP1zrtKsSSsxXgnSTx3gtD3+peXH3MEaC19r996ancUf5bdM7mYNSC/DSxNNb7O
sc1Bq6v/Ofgm+s3qTz4NReAqeaaliUnOjIFtSuWD9ySfdJmPheyu5SD1m6dfD9eLfFL6GdnjH73c
4CxyR5gLyPkw00qEQh4FOm4nskHGcHItHnYN9WEhDOYUUiOhnJggsi7mjARKtIpDLVKSZqlJFGbD
0QjSTRlsgyjNFmSmLu7u1StSF4UZLctOGQ6w2cXYT31EPwl+mVkHe9HU/5hUMxgbV1RJ5g28QZKE
QWWigRwillWI/9B5zInr2N1mmhpqvYyMWRSSNG39vAx7YVbL71mXz1UbeZ0DrjM1hLQ5AbLwDeKw
50uslofvjhjwzVwkx1wcu1w6qi2j1kLNGWrCHO3KeiXZaYRnEVWS2SX7yC7v2hW2AqtWH/pEFTmO
jKx3k36Ug2CY+JfZLVIf/79gdkh+KRtVGXstPq0/OFHFxI0DaDbdVbuITMPJhiXa/VM8irtHMyJj
4YUjAjCprSGKfFwdaveP83DwEkf04dXOMMUkRaQk1H3mUZW4CyE5wTRNKWUYQ0n80QyJ6eXcTCoo
WOABDDBFn+4vsrR1ZP7F1LKoa2v7lVRmGZtP06bM85TtQxiyLGgbRAgBwYiuVTDxTcDP7kGE+Drq
miqSiayhQAo0Ws1ezbSeZA91kYLsbhtMTzsfUUlDutB3G0roETqdiEG4XH5av0UsKySsgTrM71cq
VgerLCHC7Ik9aQ4l7TUrVcxtYRLbHugUgSdA9COf48ruFFKS+DkYPLWZgiDAiXcjKZB9h+zvGQsj
CLEm4PxYS5crpQseIjLneFFCl+l4oMMdL2fref4vSaTEJYrE2nPcHgkmZmEWTlB+3nWgoQJPOxSz
+TAzsFu2E4ucUssJWf/jYQAF9dMNMUcDmXcO/x5y5GxBWDFYw09t2Mmn0LIKFwrFwHYF8dLpq0Sw
RCy5H8FDlNIxX5WlkSdEltYG9FHMix/K4EWofb832uqMdjziPOoM2E3v51yFCWJ/lkwL807/EIh7
+LiL1cEgJMK8X3U+L+xI3tZphMHMe7Jpdht9BwAIw828+F8EbKkwmbN/3wIM1ADUcgSyKqNEe7/Z
bQ01VzvdNVTizyCb3RpGu4W80XF9UBzObfJRP0LXmhh2hyPJw+lJmeutnYvBOgHdXd5BXc+ktqoo
+xXZ2R576BW4CqAt8uOcf564ENusVpFkDeYSdKCpdyjuA4k5qsXMMw2RMxQMeZYjJiyG4hWHVMiz
eu1kS0F55lahdMSdSkqinNMgq0WKEAWRgEB2IkukDY+XoKD9g9sqI85vVCscMfpJjWMzDhn2uDH6
cs2IqkGNhQKPhp5bVl4zRrrM5jHIeyJtxy7iSq3GWQC7GG7R9fni47XkgDr0eB8Q/4DbmTl/p1ev
MXAs8TzhjYaggPonzKyihGQFWOy5mRQaxJtrxqzK99+PBrjSE1PWf+e2SNyS9iQUiRz5xFL1M9CX
Dxry3/+vMiNA9/p25lw7ZCBDfdM75Fg8ayhzH+2q5XTlN/JyFTW2VnrZEB1GjzLZgrWHJJp2i6+Y
zLO787aCFrwj8Ur0IkfgLvXHSrHj2fobLJgFbpnETffqgXoR6g7fauW3FugbaMDK3kMtsEBMZPOW
DCUPyhTBVspLHYL9Sb4TL+DDztx0O2A/1NQwLBdDPcR7wSRxs/aWxkEoIUIKOICN77wlnLFi1xh7
7NPmYX++szeFd7/pNBlRO9q76o4cmfzDVlKeLWg42YgK/CEJFfpcjU2X3hcMR10rkOtb6tA/fdZB
5plvzinGrsoUCm8Al67SGQIokmp7o1DHVSzNinqammbx0OHAoDoMacG01VJl3GtvKKByu56L0NmZ
Lp+J4DV5bUEp02HPIhtzh57eDNJnc6t0iL5tmPYacWnYfLbNQtzdvsZinytvWlAcpHmLTfO6cUfu
88VqQwPusIlsmauODjfq+5EgxkhPvr+6a3F0GRqaA4sguP/9JrIu40OfVlEly+6J3jr6Qibz1xg4
K6f3K57CSEb8VKOfS91e7sEAQX5IzeyEje8TIv8FKKSmMk9vqTzaFhoQBmVmOnKbg9yOjp+aDL4n
JDXok2HO/0+XOdBUYEMlln/24nktSaNUP1pj1bbdhA70j6qIBScCCMMZ+20KGPBwOQss2Ch4HCeG
FRKwg3A8qZ+/yu6fDRzw95XKRfTgt1o2NM8prsNZc/HFPUS9QshPnXn/YC8uxIbZw0FTwhMrK9Nd
REi5YrL3CAr5TArrwp6A4dnK3IDBFtUctconLLrI9TpwJMoP1hCMl0ltPCA2ZgHL/YzGKOscEMUx
6lM6oo/c3ba9itfkom+ZDK5EldO2eT9nMIBe7ffrf96wetPPkMkeVkVAGaaxw8mWX+72TsIxd7hl
evYgVd1/QDk3YI708oSO94TmiOJEu4f+b9xf/8gpGoJZEvp4TB8QlINeRTgdaET/gTASEx72HgBN
z0S7QgtiDKdoZJ2f61wCeFQfs9abr1HWqI31skNhD9Oi7+sMnVZwKw/KI0BtaZhdWBvc3gRi043T
H/yJCnZkwq9UMyB7CsfkzQU0GTDUHT1WYbzHpLO1mMYMykUuCyOW/lX/yUwyLVCAiFv5dg9f3zI5
dUk8Bxmcd81RRIkRy1zs0ymCUXg4dogGMTpjPsNSSidFAQU7GdQA+58rQ8oI7hY4QBoE+AqU1t86
JgtGtXShqXWH+1tnFnDjmeUZXVizpY1rJHbRhzhJ68XGNcN1JQ3iUVOYjXDdq/QME66Ewy4hz+gb
RCYhXulmakTrZpZh63cYEk4X5J1T8PIHqVKdt3uSAf2MXMqUvf7eKyiJbrDyr/jPY2iq2PJKVbP/
0GEmHDxUI4BiQevV7fbu4hmGFPYqJ0fR5ZWa3R8suvffLF1OFzN1JHvJEPOVHhYpKB05TRjQkMgt
T11OBqRgzb3AVXbNJHlidlFuH4POg3ZdHzZawLMQuNN5NjSvEejpSuW9onQIKEodOWUjlxwfCYfv
ZA3b+1i6GcP3zSj5N5KAYIrckvjWJ1wQ4I6wCBu5iy5BiqNGtYRdB0s2R0F31m4e71fScX6TB923
n/X/gIhSbnTAVoQEdTPzUE1+3acYtw0bsXaW5JUfcomg44cocp4oTlwmkiRCFZD3VF2SihjwyQP5
6Vp7lcFY8p8wz8zGZWlCOmJriCCYNEnj8WdX/6NxfIkl5/NL0QG4utrtKmbA8XZP9mxyqXToi+Ym
TTCoRIr/kljaz5UoMJNt/opoIF/SXRnKNdEW+ei0Ww/sHCOpcUa6kgLpcAfqDajZ+E2nXZsucU+Y
Wh0Cr4EM8BAxm7roEKQXxtg5wWtwO8BdsBNZ3p6E03T2mMKGOzgVpa238n5E0/hcsMrrI8Gfu2bx
Lct9bbj3fxBQPJuaZk0QZpgU+v5loR5eD6v4Bkct12iPwmse4iJ8hSA2THMS5iE74ADsgjWAecuq
c017uhBouzl1kz2uUOV+9+2k8ZmQPE9YW+ET6A6tjh2ssSA6fHNGQArwQ9QPmsJz6ZdqME4XChuC
qmFK9F8OaxLD5bh+5CJR87jun2vO0kWxndVEWdGXwd/iEzbpvLvpv8an8JwQCWebf9s+9EXixJro
8fJPffq4D97DqQxXeyAQbRJy54LoMZWIohDk4+j71mAgaJwzog9Y3wr/OIanc5G7e0bExT+q32wR
IvNBQGmjEYfUcrKJleF72Ti+XapxL+Q25JmfxFe34D31dYDTfIHH0EISXwUI/di+eEBrOdHTvab5
CqU58ZftYNdlgLObHoXHtfui72FmJEInYsNYy7bFR77MAanKcnwgaBILigqNms2r6u1yE8pP7pqV
suS/vKOVbe7dhTdOajn9qbNsp4qtcyO+tZMj6STz+om90Ji+EzBcEalk/cJ6yUXYxY41DLjJOctY
YTurQLEnU6cs98uNMDxAs2jchuupywUPT1PZpJ/Je+EC+jjx76CuMiDmLKB/y4zPrnC+IDG2csLX
86tDxJc2vZDua7LvHQCrjel76yI6wxtgNW4sgRdhp3QXzcJ2f6uyu/2f9epxuCPUwDSsKRNUVQoq
x1W4At5qXuVGGNpyyS6mdxutNid7MRzcD2DrSU1FwZNhLniOeYEKNkl0Yb8bDrHMyRyBXQS53zmN
Do/RrBoeh7tYEb7715V/CdwdOmCCjuJV+G4ELLX7o6h3WmALraxOe/laCjrcuAP/+RPvvQhCv0rG
RAcEnSEF10fT7jCDLiOOHWDqyXT9cMlPiW4+TcyDvqGdc1z2MhOMtvo3D+hpo9nfTfUL7JdoyqZz
nOiOFlPSJMoaqCECugRq733sWE1hh4qhq+eE3Oi7xb478NDF8Rtf5GBadze7A7BIGV0AsHYkNI3j
i9Df6Ck6PmdMBUCwKE3dpWoLQkV4ARcZhJDjZT53hNQuolS3yfz1Ge+dzgFBodzxtFhCbosUcNuH
epLiFY/OhCV2O7KTkQ5DYFeyzcUNIjpyosxaOc4MoS76yViFLmxHZ7xLB7+DepKyYv3SIqzE1BNr
lMujm9bA4wE5oaYmp3NMViEnIWfwbboSHr4GORARWAWjJ25/UPNxkQdY5NRjpCUjqsNsEKTW4zfA
Otkm1ipDCl0kS2oQmr2NL8dLxIrtQ0Jag6Nwu15k2qOLvgLVXrMFtMMgYFYfFaczzDSPakvXbejq
omuY8Hitolt10PCMV2f0lUaJRD2qfQVa6bNPs8V98/jO0Zt4hedSPMchisF1VYuuSXFf8Coa0z4j
1SLoI2NV+0Q4XM5FmAHaPTIstE+tcVfyhXsvI9aNY7g7/i6jiWTICzrEFqOQswq2MjBNtccMBf+I
zSB/tQp5DCNblpIuwYQ6AGHhuQXvjYSvoMMwzqBopbEPvpFZlzvNHRu/SD5mWR3IBA6DZ9/HiP9g
IpTT/lR23T20oPK82jy1Mqd9BElMdq61rBIjZYIi9sdqoro1dRtutdeH+dqZLHtriPlWWVXf3ZPb
b2sXyZQeV7ueRifskfpXNL+lyOAPabwYD8zgbM4vFnSA9m3RNeUOc3RUQyGtfq2WYo5HmfbEJXoO
Miw2E+hx8aWVqy2GTvgPFA9oxv+LjS9mKoxBvaimtT5w7aLIOtsIKchAfPCCqSGPVntArq/p+vGA
y0iMB0/z9VXlwf23g4gI1/58n8YcSavRr15K5hdsftmE4crYQRScJ6Mfyslzg9Ddev6g9YXNro9/
UUOUckkMNVmTKojl4rr0194sr4T7w17cxu3EzAZKAnJw3sR3V2CUGBi56tB2m+srGuc+110sGcur
vcJ/UxAgsNEoIGlPDZ5IwvOO1uksDAc9Iz/f5pK+yLqn7ubIVYpGKfNp6AnyMh0morzNxhicOpAn
Qgtn1OIqoXFZdkpTK75/at1Hl27BD4+aWKa/xLog7ezUZV2k8Pstzg0PtC48IrLwsmZ4Lm8ZvpZX
C4NgvPHkGhrqwzRa2yKDwRYtMXv1qXyi0SYzf4pa71HY5W5uCpjIf58DhLdPWSe/nP8cMnm/BBZZ
8tI4mrgJP52PeYlr+CSbuPCzYkppeZWZxEPhN0qW0U/HUBm6DB9jzKwX8Kx7sk6o8aiU9skWXsGe
sIbwfwcmgI3s+SV+hba7NYdAZJnOHSrXPeMCwsg3AQ216ZxYTBJMsaCmvqW2zSEvNxenu7sNsq7D
zWjDrK5HgQHcjPijzhesVOV6r6PR+ZfGbm1HxR0FjRdsjOul0qsNvGPJBLf6LjS0g1jBk9vE5qtD
Y2S7IdAelcZRfMTLY0q9fZ7QZkJ5LgkBfz9azcq5lCc2zH/cmhRbvbg/NeiPB+h+BgqyAufJX9qk
segaA8AEixTOpEzIkA/GVovzduTE1qRsg+eY2oz/mtYqQYuRajotU99x+dfdaOo1LWOrX481425E
0umVj061slzQ8cT7beiRTsYS1RR2LG5NNKn8hV/c47H3eIk2rBzI3XRcVISkIZMG8YeFjvvzwTtn
IDujOmWkOavMoToTX0N8yrkYFATe+kjVTJUE5LtltZfUMcRi7govrI8IlBeBwXvhzoCbxELOf/IK
lJgddVrS/+NTg9LD1pNha2XOe1WCYD6VLeW7+tCM4Ju0luhNkIk5vAZpW7BnHVFsopjofVT8SUhx
u9Zk7IgoGu4h4t7mGhbpqM3/YonT1SpJjbG+G4EPf84K0kDxClfZkKNwGBxJsjTVXYZEXwuG7DYa
beA9ecvh1Qg+/9OxqHIwlD21X3GUA0JQzuSYXs3ZXCldMdoZ0r8TDn+wdsPZVchPzJA92+TmLJtE
g+JCZYAnwmERn+2sOn/zJeWvmyLgfS/WMLFtDselbhOSDDCsHpzJEYvlEPH8073ItFHPHaluPILP
Qmox+dHASl9CSZs2HbwqQQ3qs5euHZVtwWCiIHQBiFa7DZY50F7MPknCg7fl0QVX9vgbveH7kgUM
wSG6zrOlBR9CsQQsu5waf8E+ZMTDdZZVVg1zBp9qipaaPGpRE6TCKnVLFcmYb0SbEOIeQgwiTo8v
hHjlS2vJyIRlNK10fr8C2KZuOUjHbUw9tsUCXQc6c6a1HJGHkkQofjTA81oulkeapEHToYuDax2n
U6xonUFZkHHi5S9sxy2N45cm1RV5EKUSW6XhtaEZchvoxVSk+tV+0nuNNLC5aiVmE+AQnRGBeibC
Di73cH+FM13512jr2mXAR54wtw9zfl3A6gpqJuUSVgP9eNX/g3S4mULBorrsfPF/cBI5KTs/ba8A
2N/AcHLOGAqNdqQw5Mq4QJnQKrb8j/kZxPOSllrUsjyIwpAg8xyUHJbsEeBcymBMUW2ihJ9SAWow
sJtP09STNKKLz87k8BJgVucFIr3nVJvzUM/tLmBlJN/n4gNryuk6OySFvwdG5wY3i0Tnyt8bmgLj
m1J9mB3A2Y0/VxW/iWJ24jYT+gSMz4dXc2ZmhUYTmvflfOy31ODOeVguv8H9T4pr4n/cnorBkucH
Dslw4KbKthphYF9LqkAVU31cOdQHBV++vskG3OYPoY9w5iMafgvZSlrRGfxknRfyPI0Lu37J3u6i
z+WNglQVDQjekigDoIYx3oIJs87vzIZEAOAbYYwjHpGqrrFxNW/EFZXQmh+0jVeFkCFS57Dpl+TW
AdpzDRdefH3/+VM7EpnHT9A6onFbGguO/hIhKQzuNY9wkNFXgLxPrwR/+LgI85+EQHrh/tA8QYAE
mCeultB8Ip+J7o8vO3cLBFJyfU3odeQ9RcpK3hthD1p+BRjSVbtp8tphLEvVPshwc62fqniN+8hl
kT6D8PBSzbyo36lOKOrq9hKQpqBWtIyoJf8QkbBMQx5+o+ozbSswShObcjRTJpDCSJJZpb/sY2Fq
PYPWRoERe4gsBqdgNEGhrfwRpqKYRefHEFCEMug06Z9RKlr5wQ8fvps2RlVmeZ/hLpruhJkSVV9v
sJq8FpUXwsnEjcEAoAso2AWCP0SO38REyYJY/GZ9ahcIBjdB0/x/d/ZQzXq0AFiw9jxRu+0Gapgn
bIVi9AJNl5ae9aWAwgij7U9qRHLAm5zTMW+cd13gUjaT/WQPJ/fSl9IOkY85/ZPAcGVvvMLCRZ5F
WBowsGSXVr2ESDeNSvlj7G3PcAZ4tQcUXUDxPnjRJnKDBtYTiG3l1rwSI1+hUAoH3wWW1jx6ygnk
kBI/l91r2/V8NZf+/UHwSkDigu5Fplq5PeCL4fCJqG3wkd5Qv74PDt6f3GtLBmJrrzCO80rMPN3v
M1WQct7uro6D9typ7ctbaqqj3yZcf0Z/uIsyJu9alfxioKTcgo4Q8P3oG1Rg7n+9RaXrMNnLilaU
aDbYtpaGLkF/rQiPVHd2GCUbr+XN68QTKXEPLJORCGIOOhDcjKXn0CnlDD6RG3DkGL0j9iBDjW48
jWLpp+aTY5ttdRa2QOGbVNWk79sx/u6bBKqdftoBrTwrDzo5OmsgRBvOgtF5LJijKHAO0L4FQTHI
L+Q5e1NY9pIpBwsumfZIGjYXgxyD32P9H7neMI4JVbFS0VBoY+fEY9SG85xXdw27XznkjoafqD6u
I0Y3mTxZP+NOt6qTp7UrSwVsLkLrHsBVWEAkZLbQgcNGOFsPzx6IBOggUVca1cOavzsrV1KJqe8F
kTe1M15LbGFp7B3uQm5tBW5qVREOYUh1RIn5Q57XkQI3Kv2Gn9c+Xu4RorX5/Zh6BMgX2c7FzmR8
W6QDXqqrSK3OcH0R9oGsnNhb6OiQHu0FPLro9GIadWjORYlvqpB1PRIAZGShetl+d4a0Kpdioq1/
m9hjisLq4HuIeV/UDkSGH3Qu1cwZsRyw0q1tq9jTmnjxGZ4Klf6JE5G8UlCmf/NJanSLgnY1DUYm
rdNu0rO9GLiL49+uyHPRA3NAW7sLGMbQNnz4IArgmZUSxGqQpFWgc2kxfFXMHirCx+MrKdCaB8I2
yyKWYvWX7R9VlZzWxs3OEhXkVpRkXWsP8YY0tgzFT2q2Qym+Ajt+7NSNbciZ9XdEOTTKnXFVBldS
IrPHNqGa2iUsmKLoj9Al1gZhjvrhOZJfmDoTcrmlFC3W5FJuJx2OE3xOxLGJS5Trs1SAOXxIl1Kt
bTZnC3moY24Ja8oCbDm9GHtW0rao4/tbVXSF/prgN/RHksAJHk+073avpytfe75JmvVdWxSuTyer
SGxVqc8XBzuy9ppr3veiQhAfYfy4KQ6m3IkFm8CHTRlWsHbtKdfhmD7NbL/0H7mAsMZwiyQvHpmq
bLyHi09ack0ABZtsYPkNjtPUI6LLQiCYn+DB6xYcZ5iKJRTasgAGSsk5HiaJjqhkKu15sYkCX/hG
KfJfyfdHj8Ms+MRgAvSAWwGpsupvC4gUbU8B0s50sE+DnHJiA0GASzC+HqTPDT2dkzR+HUcDBo1w
xvpKm2B1GZWFmwss9RrvNQyWdJu1VSkVMfX77QIqIIUFOvWT9M/DLWzuVdwTYqCkMo01inom4hEL
5W5tct0q6ZNHP4XOaXbMhqxVwWIzT+EQs65rYxco8eEJJ28miGKgBypWrz2oJAbRVWk/fh/lM4+K
dB1OSC6J6cJ2jSF4yCOkzxJwdc9ztRNI0qZbDjiJxVp8f2cUst3OM1CpeRBoJDp9glGpX9sTavHH
tTXcJmqiwFvYINJ7o6PKvurON10maXEPX8Fk/uO5ZfhPCJuRINFu0QryPML4LtmKAw0mqJhPHyVV
OmJ5WcOmTAaWpXG57XC96fyA2OrFpcxN70b6tVLmgiggU1omZeBDjakXZevjnlu1pGhcGS7FCSlU
6rzVn5Nwpypk4AKPbuDZzpNIHecu6WUBx61tb52zRDFtp5L6viNcVwQEHJ8jhaDl/0dFMppeV3uV
hTSRLBCBs7o1Z99MWNYntvIJBqpyKNm+v41kPGqvgFQ+lIZC6Kx/WbVZt4I2dDuYL5oeIeC7oKRz
Zmb1B29gv5EEThQRTxVdAJkSc+DA4dhSlfDG22ip1M/reAsSrVHb5u/XF/cHqEK/4V3vkU3+HmDw
NIacRB2I9staP5hxnRb3BwaQy7WEdVSeL91DbrD57K6XJ1WKpAKmA7cHcYHbc9RA1qsnGRvzEijl
7SMHw6HYeXaNd5Ww8tTSdkHcFTyIkBJEzi9CptxvvvLw/YTQ6MeGVJ3UfWu/7v/zyGUwPZPLCbuy
krZp5lASNyGyW1emrYuwgDHgWkIXp+4OcKhfuur4t4XRtE7RWYHKF0HI69PdaANDUKhyNy6NkhpX
v1ObAvIm2gEiKFty8GCbNTyiVF/Jiplhbw9lg1jS0lfisdgwaHNwOJ1uM/TvwEzu7MckBXPwlaeh
O4BBfQ21uRxPSB1tt2X/FluJ5AAVMu7I/CZDpwEgUZ7fApDkZey5LbNHJuPW22xoYonwg90kTUXz
2tBHD/w5V9XuKdsEsHNv7aqTn5DMlmhXuybri8dfvWUBs1aGX02159z/He2iTvb/GZAITbelWFaD
2UGw2dLCWAApUMLX4o8RF+fCSK9nP1QQa+D2eQdThDeyvAizQ3mt5rW0GoZwBdASN7Yr5RyajpYs
i5BirxJ+27XqMNvUnUODK4F5Ko4V+/gFDC0HF0x2GjDbMH0LRlAL9lqA/CH65fJ4rEmJDfgWgcp2
VjztfgJJDBKCBPqoB6dtfi6YNO/3EC1SFN+s6aJhqM0IAutL8+indHD/E4BaJWZh+DemxRY4PlUo
cqGc62LMtyWrpCy5fu970Y2T1ccSUxY0bKd/9U5AB8anU4AJMIZ/F4dC7++uybp9dJaK4klxMjGC
KbVHoOoF+EgOlhffUsdT70dFKPQQHKslV3XYvFoyYuRzqlAFZKFwpsAeAlY7DQt9soIdSf6ed5dk
wEwVmFMtULTfO3V9lKyFn+i0psnD4THurnWrCPFIfAb/6UZ/jGM61qG0j86AKQHl3GF3oGovaaOB
Dy8uQta4XNWNloi+s8X/Gzc2K7p6iMql+qZwZ1q0pbLwGQR39g2/fzt+JbwXGhteQXNhXxS9jmsi
0jgC55HgvLpnnXJAO32IEyN1aph82paKvr1roypAQUtTaG40YHwktowSX3aHJRmVTLYlD522BOOq
f0r1tZlDGYNxkHkIf7caq7eCLiBYPsDBKWlvV+8Sb0k0FCcyUmoTgeUNQRtCZEFsNZgjP9E+YdCh
ySPhnWBjQWVvGfjufOOBTSgxKtrOcz7ntWoWpZdxLUBDjNROpyeF2rvTRC5k2RlP34fYTJEWHADP
41LJT+4GayAKWcFB33joJMtTPjm6FNibNv00QJGTn/OR8fto1J0itfsU439hLwu3jJKgRkKqVPJv
0hrM7IU+Zy32lMlNQSrPfZa9EkqO447Tv8kd+tqnIy6xAp0m4Acs7bgIZdbSvXrWaWyOA0FtRfis
9CArp8pCHprSg1hg0JYZPfhgBFvqg9gF6GyELRP/wke7sP6p98QLtX4oKrGDuqAP4j/h0uCEz/mS
fH44si1h1xVeROpIpgmOT9mJwYBajFa1wZiJQlZU7rcCTJfufG29ZgME9Nq9adKQCpHueTnz7YAH
hIlVPZSCYvPRFgo+4uMZYUJlcFbUZ2b+oMz/H18PpWkgUTjb+F1A2fL7Y0G1k4DWoQ9oGKSOKOs6
zNjDPqfg5V0mXMoDV1LxvuZsw2WWIE08HoDsY/I49NS+rz3DgzuTvjCP5EminCaKfKSoYFKYRXT0
hJYYL+LknmVOF9//vylkTxEdvImjjk0dZ4Qdc0hBIlgLj9VzN4AU5CjVGe2cuF+08LmXY+bVtgUA
XyhQWS44I+KL8NLRRFpW1dgj3a4F0YixDbXbTgS3T296HDvr/ZdrXNA1JD+Kn68JDHhjqEliS3Pg
Vs9iK+AaBMMkUp1+WuYMK2eXJuVhmH6GH3IIAkzHozgn+2YkaXJHOZdNNnFI4PYpJAxLUEiKoHr2
lXiDKDhyDCZL889mGVJDonTxBbdXvdaOK+blZBrF9ZW1bDNfpnh1otX4PGhBuZ09S0RX4BLRcCQH
/XOcxqT5bjruquoVmknvqDGVFCt52dHb4XN72aM7ow7411qZooCRoUP9IzUq8A+Ad9RIxy4vIku5
6eVKK37sWhmSJW3wHb+Si54cR1YPL43q7rtIlVOwQv/u4ULEwMy0dEHfkum8aqlx6ggOQtzS6d6N
SHlb3jDkg/jULnheEUvy6UzibIxu2r+gV6BTWKtcpM999GEzaa5t5lhCAQsG7aqV62S/XPfX2uvW
5yrpAOxp3iZAQGMXro720uzYvF6DFCL15Vr8TqvNtuWX+SDd8N6B7uXf9Djnv2FsZpJfx7C7sWOk
BjgUTW20wyRTjHHM0/6/WZ1WkROZWhmvko6arghuEPmdEuT23pT8guXD3CHIFDPW0Sz2dKvh6prF
aR0JBVa8efen3Oh5i9F+x8JtYDbBWwEeq5DWp+cc2Vx+SM9pwV8TfKWBRsx47SmvjMCqBYEKwcKW
VsHicqlCfSoz8qdcG/NHtmN1QMdeA6TemsQ4aiGQ1z4I794KC15uQtxBXEtFCDvxd3Kyp/1Nfn8x
1LQnzaZ/iyp/Qt7XXgrsMcnNf7bMnlu+a/A2nPk6ThCMJHYfna3MlmIlxe2prK80X7k099kmnotD
acoG8tgbP/bMzy3NrGJJs4DyIPr1JYoXKhv5Fgze7lkRSVL4mYqAo8eIcZmcl5NdkRFLdXOvWqIk
0+++qkDk7vxKw1l4uP9fiZ8A2NqAp5iupfi+IK4lCJ5fwVswAuDms0vWWxaq3pG+ODBILkeiqfUO
NxvndyZuMuciHbkWCxQwZaWOoGHBmj2LhCJPM9C2ir2KAOCGIYHyaBZR4P83Hnqo45nwnxcLHPmP
VXvEqdSw8+aanCTJLXEbYo52xZSvjL0paqzFm/ZG52FR/A+Nlgt3j2wbQay3jFDL/wZb9pEoZvw6
BJhCb5nap4fLiexkdxH/EkO+Qk6MNAZOdDcyFO5Txf3g2Slczhi9KkHkVDWhvWmMxgz9QBZm/33o
QalwbDoBC7ZceZskZEiQjpX+atYVwjt4Axtmy1c2iUdhkia+vdmD2j7ad83GD/apMbyMkEBlIISf
WpRgrPTnT2LTZmDxy4lgiWWwlzkRFqJy61zXnyOt4yIdDSCyZo6iu5XdtA6A2zTlnQrpcJzc6+DC
hsg4mgrasR/SNe7hV4hqyeA+XlEw3JYr5t1pLG/VU9KOJRj6J1RVBzgbcPOThzvLfeJcIl01Yol/
bMkolFN3ph0RbaAl40EOvsLPFn8g+Ng5Kmuw9KW+nvW+taKTOYNLVXx+9D+TI+C/9jI+HSMXeYQV
5W9IITtPQsQHSrzv9d2wIVX7MNsAcBDaYBaQbG93fyrFpUAf6+V0uFPV+KOWzNQuSYreqJVydap0
JgEa33Iz1m3pdrc5wdx+K3g0Lqys4V6kbNOnEqki+PJYjT0h73AH2Iu0iG0tracJ8izLc95zzYXd
A5SgHLQJVHnaDlft3Aw/MqvvJSUBXcY5mapu/DE6BrDVCORisC6Z1NuYZ7du9vn1P0j3yg4FW3lZ
kzYJMfB8owUYmrR56VcbdzIthJAYzSXoOkFy5PM9y+hVXxFCPJDj0rzT1rIWRQjUlNWWVy5kjlhf
NmKxBXlf2iE1w2MIx6aON5u6sgmtYOGnQbtGZ7SMSvRv1z4/pa5dpQgT5JPy4O5jPCjlduQ2UMxz
2/fw5UZD/v/pWQuBvxrnVyubeqBm9kjJNPzBD/UrnIHImA42jb4JWVMuI8uqWhFazXkZtQUESaaS
2cgv7hIA9Tz6tTSdX1uJGPk6H0l8g89b06MD5ok1TqHOe7atimy5i+C8sDzLL1bQQzbeqv9YoZdK
76CgTEYuIxNuV+HligOrNACG+XaXePfTIuSHNjiOmAyCyYzsH/iGJHDZ/pPu4fOdE5Scqo6VEv4n
sHAmvcIAsl7CfdYtGlPCbeVQZAvOA6EYrXu0uvMv8yxdKlBB3aeW5O2QbylL+2vbvYsGH2bhic94
UArQT9JW7kEY3oPOhWDFprrLh5GTAbjdwXfhkdOTLwgJvl1avkhQNealpiskd0NpS0Z1us46Hq/X
ezxQSlI7KI47ok89yah46e769Jb4uM3Pntggmt8Z7rC+6h5g7tlK5yeO/XSSlbQjeBH8Hy5w5nV8
vrAZX0yvU6wC8Kfrwh1YzhVoTpB4kMEitXjwi80BFYOtATBFPSsNKkqd9RFNve0CBQdiUrE+Trau
Pd7ONrA7EtpkLxpN0FK+j0uEOqzbDq8buakwXm191cajyFhkpw0y04icYEN3C5jhuXUDfkIHeCU7
/TlC8QdDEUL2MS1BshKDIHcRk8V8Ie3Z5uPI9qqMwTeX0tY1+AyjYAh92xrb6LCgTH8azxNA27xp
k3a3iB9QpEBy1rLNBlFS6qZX9MarplkisHV7N2foKK/ljRiLTUl3wqV78FOL6K1E2/ZgGrQRVRyC
lDfQw4uedR/7Exgfvy+qvqkjFbwxt6FnxhmyANp1k/9ksTG+5rGlmlG2VbK3V6d7+fyTH1pU7QnG
HGqr9xCUg0wTNpNUF62SV15TZQRNNJtbJ9vk0u2VPeBN6rMM3zpOWO8/wY6Q2SxS3Ry0YDLpBgyy
EKOEf7ur5vx9pxLaPc6VmWsp4JKPiqIh/VssSrq8xVHKPTZvV13bzHCgc3o2aQFK83a1N/V11nhz
HrNYEfmKQQOWa6dgPi+req1NS/3mspkVeT2OyJOwon21rnFc+iUExF0QfvKnnPxQvdVw+DQ9swlJ
Z0pn0fEqg//4+q9D1aCPDv+0hIboEL2NqdL/69EHbWXfx+6echqircH9CYWGPF308pCW2pX99+bL
/cM/eg6wxB6mKyhJCYP5+Px+aJVz2Zi6r+oUCb3UUklpKtf/IcUXoGpZAuWSVnrmXPXXAMkA1Tn6
iIYCi+ysA30VyCVdUPheB6Cabi6PaqnJEHSaTOwe/GNMP3M4HfdVJKymnwg/Kp/Z9iHOSBIBP7KX
Z5Yg9xECJz7mA1YY1H2X1bfJAJSEP704MVG1s7K17psIuF9uRt3Jg9q4+RfOSSAxgaIEOvFOpsDC
VdDojt3IEyxaHPBLNjrrR6mI9Q70xdK2X0Fs8tyg1Jxa2rXe01vx4CRy27+JoCIHIxEj1MdakFjQ
bN6/+4pBkwhHtaU+yLtLh3MvYqYqKK5nDzRB0ZmkNjbEzwWd+Q3t8bhGlXHxamNGlNyR3fPQIseH
lSjjUCeLh/6LGkH28IEFAitCryP8qsdD31DDPEIcHGHFUJ8BcVeDbc44ND7PEhVy/WSg16RTshoY
0xIfb/JqO0++C681aPgObXqEzQRqWC1NO5DBCKAcPl2v2iZqCmQ0fLYtAYnnFn7ixkOkxMuX2nnI
NXYW4rRIQyG4L4IKsJ1YUU0aDnV/xXdwXni/S5pTEyqPyEGX7Y6NvvNq0G87HTzS2A2kVpbz1Amn
CwxE+AXd4QZZd79l0mMv98Kaz0tNPFq8rN6v5JY93faKJF2BmiMic99Lm4vurASrqwy6EwjTA1vh
eWZG5/BkKMSuM/zJ8LLnKcVuUrRViS53BPFQEMW7xrtdSD3Hl+k4ZO6BN+j7rjrU2ZNI8nnoRaPP
1meeXuwe22L0qmezU+rvhm24wyRl6mGxxXWD8pNs5TYY0IpaPdUhKv6KPGA3/B9XP89d2osUKGuq
1AZZBoRJVhl4qvDPU6pAI8kjjz1FTOGayRAZJacpstrekjYkGrBD/tLQKZtFsd8S892WQofzcriK
50qx0u1rOQ70yC9sA/uZW0S/b56CoGBDn9aDe1S0m+E/WIrE4lhR/Hbn/WKZp43iXNoLqzZ+7Vst
Ayfny22UHIyNps+fsai6LMhRtx5Zy/3cF4NCt8T7/Tu5jpDVits7cWnQfgJlZ/5aeUtqzzbpdHf6
OtBaLNTJomZ3o5pGjQTGsfOBENK5AVYSS+SsV+/GmOhP1lJrI3o7fO3SVQ3F3dZUld6SZlp0bbs/
tJeB6+WD8MkvgFsSsjvUuDBQo6PFEA3MzvZa9vfRzr4U182VhGyEiuUGiHJOk885I9aomnqqx+9m
hM3JfvHpSM0jstKMN5SH5dH+wbQfYLLr0kFGrfvBwrvj8yydM4bxANCalo2vL8DbiLSRLcnsi62N
udcwFPQtxaI+z78Q9xUVh7OSw7B0M3qrQaDasYovFMlPjhVBXE/Vqh9wppYLMqYobW4KjejEsexN
tTZv1gpJJaGhvm91U2x/oCUNa3BiKXEuBvMUwSZpiHFK1Px6J6fobQw5KgKcZPePAsZCd9qwF+g9
4r+5Uk9zTvUiqSG5CEAPcAH8NkRBx/1gBs08Fh/MlkDS3H7GE0hh1Dtylm4cfxDOc3CVAxEZBZWb
kyO7Ve6hzy6lvFEalr/cW1dPAG1UF9HH7+eed+ELmVMdgQeb4kDyxfoiEUnCTT56rlq8xwVDxSVT
ugREAhh0879+bP2lLME332qDG8lfVWFHqufGlFArfv/JPEmS0rESVVhiOULWZhoIKjSODvqnE1Jz
AjvSnLNilxslKt2FFt7TgdW1YB+mHClPPNrm8WCqGMszas1hIq/sXTHc6PDc0VcnBH6J2S9q8K8I
fyqhNQS7IGzVHYzbsgQY40zq5N1jzSQMffFXj/SpSGyUPo2zdCxoEF3LdC0KcY9vddrWKzBscuFY
DOIXXYiwASWltyYqdWGo+m+0+gQZFc3uHaVstIINqRh+TmZQKN2OUaYN6OGYcl7TMvvFstMiHvIb
RsI8t9JPIIID+P3hsln/E3/Ykvy9CuQ+NjUYhdi+0pmyaoI6hb2zaZVNXVQmyyX4YYBRea5ioH14
T1BUD+j20Sg6FwwgbnLPkPEcJXbyWiHQQRaBystWXy9WdP5JBnic/QVZ54qDhED2ioEBrUMXNJlm
atR1ZUnF4oe8X2uu3TQ0gt/rcer8Fvc9R6FSksy44wkIZCb/O8jgjpLWae1trT/WnuYXeItAZXMD
hC7E1psAZ2dDrE62QFVrq2VxB5VB8maXwxV77QPc7yGmg25xvJISOhZnp5UXARx74Y7MBNF0O3Wg
zSliUcv8gokEwS4C0XY7YcSVOlxTQ0RD74y/MOfIriDti6Bx5ES3TUjkJ7DWso9LoxA8xfiCnLHT
dodpiyoFP4MdcIWFMCku24I52ppQYuPK5DwC61rW8HZT48Ycrl9AoIUyj3yeEozImHyaH37GsVyR
r/Vuf3Ek6einpRcBtyYQVUJTQh5dXpLW+q7eVs3hFBcRlBY7JaCnaGGr+py9/PYjMn84Alw7D+ai
Ztf1REnP0CA5ZpgDhZjCDhDYGBsYuFatF2EWQpmMxymdmL+JbqCbkdSl8BTS/wQAkPBUFjh7pUgI
5oc/1BapRRFzpY7pWxj6uFwoM5n6xRpeYLwe7N2qaxf8blecYgeb1oSkjcHw5zAJW30gVNHOscHZ
yqsYQfYMNDNsPfhpyd43Luzgz9ORwN1zUqFJgswbLhdGFjCZD28WUEG9H5WDNdvzcZ7MdX3PjpZL
ILzXHGMR9GExtoUNPRLIdYH691zFMNaQ8W6Z/j9+KWT2IuDJmTmKZ9tw3EQbMzWE5mQhmFpFvj2G
EWt2CDz6f8RrCabrUxGkxrX9vKuuqkhUI2gi7GwPozfAHlyg8zvV0ehE1QpDp4/zUXBrpCQw70RX
vnAioBocIyR1xNpv3hr6r3r04Z/zWTTdFj+iHO0g3OZlvjWQ6sN+8XjcKfmpPFUZPCqK4p756sgr
YRD0+oS7kTabw8leKthBAgJDbCR4AgoGqRmd8EknF9wUcGsLnsPDBoTgg7/6P0XKOT/Bv/nJ+f5i
PKKLIjvUy3Zc+NyUdRAZHAsyu4axf9Wl8+0LdijOL/INZ5W27+uElvLeWRdjjRO4JTeIrwGWbfBC
EvDp9wSO+LEClFDu31VQf62IORCBgyOwpDLx6bTgIlgeFDj2GRX/ySYEXq5wg6GRyCHRYLK3ClXo
OWgkE7k0fAREr/ATJkzkpn+5DHLKakBSnMf5Jpie1WvZbepDKbiFCi3+M8jSjcG/YIXnrLNVakJ/
t3XIw7vMtUGonYS1fKZtfjfAABfzVHoLnHV8dVIcR/UCxr0RFaW7GMhcJXS4EBeXhQJxbY+yiXer
LxaSDBOPMGfBsHGw0cwFzDsQBCjBIGa7OR6LpG84nIbYwsuI+Q7YUpaA9tDOMysEtsQ3k0c3dJ+n
Ys2G4hEgaj0IsE/Tz8vXZqMHq/iD08rqe7cBGYoU75YmGLkqt2H4aGCZIqfftFJG6NIf/CUpY2gZ
65eCYxWyoJyu5XPd6DNCUJK7/kft8JFzFnZY3lYcTVbZbHgdJTEOugG5kVW4piP1aP+cFB3EcoAO
QsBwbrrzuSgoQPX1FyojCyGYXty1gNf4kBtGJmyuPnjbvhVglVWFojT2ignhaVnvETIlJWsZykZx
wH7a7VNTlmOA0pc4+695m/zEI6ruaWKw+7R92Maqfxt7RFiu0UJSwOhGS15OP9A5yDKvbV0gdW5i
nxDeXRXsMb9RTJfjU6hQNgnCu7DETUZiK45E9ozHDlnLR2qeKOczkq6tz0WankDd9rShk9Xheljy
YG07ipY6V7OAaGlavI7bKoHIjXbDByl7aAWSv1M7BRqBa4TuoYYJgMQx9MuWMHhT8iRkePIIzbQG
aKhJ+16F5X7/FKJbLAwXm5fkH3PFvYmHnxrVEbLv5Hy3MHJVC6HjlgvI7iVL6uqDBmQWj01Hv/I2
JMLJEK+vYFy09eii/vm8xBnmZ99Yd6ZZQpHAoaIjidirto2KvThSDNb3HF4W7VbiL0K2EshpM/sm
STNVvz2ojSpU0aU6j95JFbpmfZeN0f0FKWpzHV2U5aFdrZD+8565jpMGkgCwKHHxcyCDutudnytr
b5h9sZ1z1EL5pVTqWeFR8L4ikIa961K7iw2Fc0nyl0LUvdCKcmPEmAhBFCC0RN2nof8KMvGp3pEY
NX3NKoik+o8F+hpJqyGsUeArdyjb8RYm7p8YN17zORV0wsnM9hR5HTrlyTrbjBRo5Uy1LVuJDr4N
VQI87euedeO59yW8cjznDveya8D8hEO8200A6K72jfcvus1yC8gAiXHhsXbz5s29NhTwxmOhfe6y
QXxSg+oWdhAKZtmkhUNqWjL53zfxstIk4YhfexUhVYLwQPSSNoV2tI491QtKDHaiwu4M6F+1weaY
QqvqG0ckKKs86JM/DHVEgdIbWTiEbNRIaum96kSptCpJwM2xyIjmz7KH7Pp0MBWygM6iHe5eDpdZ
ThfKdK6I4ep6p4T6luuWeGcxALXBtIKD5Nt2S1iGuoSSifZATqwqyQ5rhS38TW4hWs/97takKy28
LQXCGe4ttJvkjnlnDLQWWJFQeGFPSZPCiaFu35e4J1XwJJb9K6/eDY13VZtYiPEqCgs4rIcBhqsf
bgNMVH3Z5BtCIfhSt/L9tzxz/Tr7bhRIVt3sHOT21hKOwzL7H2Xdrs5Koi2XSQ+I3umtmLRw+m9G
hkP9qxJp/9f2j8Zdy/Pm05L1auWbxSvMUGAOHthuj+A0ssKG/45f9bJemstrQOraPBL5Uybg1zAQ
F198GdVk9H6bVfRZtP5Bvev0K/vKUUR1d/TREWbMcBTJZjk8sS4dWhuaoDGwpjGWtNeWCs5KyocK
/HoQZ0BNf2runxmZw/6XlViGr11/kyUjw6SEyTsr5xzXbZtpJtK+aP5/AHQjbQ37TdT5KYoO6niS
jwq85VY+mgx9X/GYW30IGvrOcxrUFnx40NsNIiL9dbnx1zlL3thEbcXdCEJrcJ4f5f9zdVS5Xx0g
iFwXy4My6XcriZRQ8Ha2rWIw32+23PONsr+tEul/A6a8CRmpD5lF229O+CwF8lBHy5jEmNiLKI07
nuGABYSENZ2Wk7lYVB7BXVdH6V5c9VpJEMXaedez8huzK3PL7W2UCYs53yi0fL33zJco8OY6KZYU
PNBDQwhJjNzqcLBm7x3ZTmIDjwuADtmnb8UqNRFilqlHUMO9zDMDur4tzLVrRWRrRuqmvjYtcrqn
XN95zKmAfavPfJOUE9I4/YPtwWn6cVXsPN/G4o/6nwG4q0kc/oW5r/ohZ7OBIIkVayonwSiLdEXi
J9IzeuAmdHGHMn/B3tBVU0apwhbRwOE6REpuN4Zl616K+RR1akQgOXlyysj9wBByavSKtIfFUmcI
fDCDCfpnD5X151Eo3uFIGokQnmmHRLA+GPgAoCGoP1lrCsMslggF+xApZjWyDJePokqN8blAucj/
o+VdgFNX0lq1GKGQqGWHX/In2kC0G03uZsm27hf5PahMgedn8vQjeDeB+3MTUNH1LnM3APLnnat7
Ltimf4C7gZxW5NmApyKoaMZHXGx6sgUk76vny28T87/2NE8TwaBkVUp1AMVEJ+vOx8qQ8kUB+IFp
0FdfuuDtMOONPo7B0gzIh+BRJD32fxxptctGc05fwICU2OZe9Bo4EKv1z46l0gRq1Xy8Zz5l03+m
aIYlQyNyRghT+Ji8S2lDXvfGJpOFJ+3ne0aeYRNOx1KG8XiC+5QTSET6q7IIRl0M6/aoTkuCHE3u
ujmVyJojapONUaECwNyvktbpCmqQ4q2IDLSGyXXdBrinKw61kBHg5L7J2BeJjlPJoRvm34jY16dX
4RswPd0Z5uGJKIYu5juddGcYgXYjzX6PXP2DliYGBNBMponulWgr56ErH17l2JCJGbsVhnpCBEhe
kJi8qjR+2afJQhwOpDtrsmZZO2DiLuDKmR2oJN3ZQyKI974b8wwAwiEvHbi1+/i04ZvPa3BKv4TP
1NpraGEpLsmAfCrEJpebH4AaEKDlwDlbgJMh2axE2O9Uw2FH1mcW3MnmXHCbgTkSt3FRX0f3bBbT
nVcizuUy6Lp268d1495E7WVqp5en/khegcDFuct5rrlwteEAbFt8+CDNQTWShluj4NCukoTKuBIZ
3U837QnUdxrSEihuLtfTQQ0yRvd98F6x+9jY9ciCYLn5fW7fbwEypSSHpBrST8lEKfNG2qTDDmK8
igylZwAvjKzWBoxh5rvaM8VGpkVaCa+TsrK2eIuHVJxritZk1u75Ph2rl/L/qXCpiZIgyaIS3LKI
vt3W/piDY/1GB/MvB1/oJj915Icy8S0fOxsqjjMWii7DubWgQe7bWXp1ZoGf+inG9Kf9xhmvWknk
HtoJG9xaQjM5FntnTF+H8vXCTZ37iqPqWVZZYB/lKj2yqHfoAU6qx4awh5DfydIrew48knVP0s2V
B+6SYhJ7CI7PXmsAqSx6NNDTJ/vnW23kD/YUUn2QX6WfGzbgenQoiDFGfDp2tgjlJQw0iUFBVAsQ
PSVtWwzuG/P6tJQBdbZ9cJSbQzEyx7szbr1DI5Ce+jgEtgLRuCAZ1rzLq+jlpRQJGstez3DMBm2I
j6apJq/+4LkCr9bhpxCrtyWJHvzhqfJKH55/hdnf+p+jU+KLND4HdFL06Fg0YRAKqWILaOWetT4y
WH7PZcyvYrn6MYMXg/wQbAYZ0IbxZEfF4bgoGqv8M9565EEoLuu4ei/7gpUUuLi3URByQioWiyzY
ReJxR1PlbDTf4KCZP7vl7k4fwZOWEHfJ2u5MX0uoVvQKTU9KwG8CvUI0duZiTuEeZ7bJyVacCGr4
o46o3g93SU1FMJGnPPLE6Ks4vjanwhz6uC0y2sVejI6yU7Y17h7Gz49FDNsRvATvrnE9vqbR1YRZ
ZFjQk/9gH7Jp8Ua52eEACGCxhysRiuKrzbMzS1KO9EI8fXp0FFC+knoGTvsVPEqnUvHV8L/mvkI3
X9KBasypK7JGCP1l0hS7lRu16Qq1ErNvfd3rtkDY+11l1f+S1Vc4IK/thq+YhGu4OVHQfgkLlUhC
pTJPc2q+VnRsEdGxV25nErBHyO10dcMukl84dAEaTNSkqxWqa0iwEvOw+7H3TVlliscVCowa0RXd
DOKlROC3OKSZOFAbbISRgPgkIzz4M1f6gInlbc1FY3vxfM95bTsvI44NSC7BmxbW3N/MulSXpawN
Ny3pi0K7jmPVKsfcQ4s0tI18BfLiVVo47+QyBFhTbQ18Qe9Fa0gau9eOWdxXOe0SsqlYaqJk5rQs
dRH5VXbXHZY1IGZgK1BtYwYJvsjzII84zAbe1b7chkLYmZ8Hj4XK0zi3hy6c7GKIE+tYkzMAYhX+
FGcQpTAOO0DZERf07QHIDV3hCt3MKQKnU8xYj+k2o4K+pFOuR2BsVRTbRDdtfDsngTqCJMSWeGHn
Iu3xbqk4loPzsLWn4Gr+5WgUJAfH43rfEsBsl8DQgJIN0ZAQEWpt81ZAgNf2YX3Wv5cX50NMyzsl
4az2mqn4Yvca6xy0DVEze04R9Hzmlis1Gf9e+rfk7x1CqATUQ9p/RyHMTJC/LmUx0k32TCx6QnA2
OMkNaEzCv7R20aNEySotWkhWT2rLKOQDoXbafdy/gS3XbM9yKiAO0ZKvkeS/FaumPB9DEf3klwj0
rRYxXxnW5MnkDAIWTAhl+/ELu7j2Uym/P1dgGGGyDK2eIuBvtkHORe4v+LzDVKji+PZTNFXLmweh
MZdzSvNPzKx4vfFuEd6SEdxVE87ktSOxUdR0GBZrYl8vG2HR2Ec3UVMmimhIn8mNNiFKoZGJlvz/
jXCTFvHbjUPN/dLw1huLjTgxmHhuBR1kCX9O6gOB28eIbGfm2pTdaetebtX1SdD1lX3vd2Px9XFS
5/q4UFUTlEFhfBp8/yiKwKd0U9IPsHV8GGRs7eMMf7MxSs0fSxJxLmQjTZxpbBZfnNPcqB0slvPE
vEzIfkUVmPNBQVaXxYQE1yDZ8Lw4woYTRybdfDKwd3UIN44nlN9jdDU/k+anyUZ4ClDIhzn330Ol
i9aHnsELv4Qycz3iR+tiIGwMHbuH9KPxjZYTFqZ0wLUKtxHgC/jNh4AaiqmuZOB/JC/5nmXU5YSt
NsgEG8CUewRFej57SHGY3r6H96avl97k3aWZudgUZSZFjwVnlabxrffglQbZhNrSOnIhRagsoWsh
GbB7ouWfl2VITqZgACWVjiGF0JOem8FKUYLsqQ+KGl4Jh/BbiLZAGPIGe+NnJoyDEAzkyX+Fh9HA
bBe4BH76UOWPfUkGcMxSrSOM4TvW4jwamsqkmmrHYNf6jOSYvITXHqaPhcIqTt5ZdQpoOC3HUvRS
OltekK1GaxizaMXfxC/FVnytvQYRT0sjKsEj3LuPmYUVEWzSuwvjYzP7XxIUfavP1WGVVPv78eky
I2K5oKdy30gvYjPnYO+MOP1n+KN3RyQGz0Dh7EtF7Xgjb94rt2vy6dkV5W7gN6Xglep0lPh2voTl
whCztTg0HhYHvY3qsB3tL6O3UfQFKmMaLb8TIEo1Bmu0x8vbXhg4MR/JSwyvJHr2fKXMmnifyJsg
LpOOD865stEDcJrHVAuMQN7GtLAgMCAc1pEj1trsDolNx982Yrt53dFI7KubpPw6WHnvBd2v9uuL
s9MC9nuFXPaT6weMZgm29o/XwK/w4Ia6boQQEi1MpIQcTQLBquTxIY8U52R892YENekuRRQKWp4k
tt2lfWrxUQnKo+Rw8AXdT8mq79FOcVglxVHCQEvknXXM6sV6oPGHWdHbV4ymbOFc26DoSYGU9U71
ZTujz+ytfpWrR8cPW+3Gg5kgROhnVoLpw9DB1SFUhNofuT00LGkIIGlWRK6oWirxgyrf8sRyJXQ0
ntoxQhQNm9cakGDCJMlXILssOHmh7avO7rq28lUYg3//7eiZxU3T6wY4gKaCOz+yOHevVa5h71ux
kvy4xUtdyTVEzwBUzlNAUJUjBLp9Wz0ldbeZ30sWQdaFLzICeD3h0AIx3IN+zMW6MsOZnZVTaYbY
e6WJaTSLk32ciGGcl5b1lYFXygHfTEYGRdk0QW+GBczMIfGb2ASZgs1Fnlj5lfEpPJVesau2LMb/
r6T4ggGzg+igSs/Su5XegyrxV2oBuF9rDVzSF1dphexoNxv9VVXEAxhQKcSrwP7uncuIj8z8EJN7
uhjEsmXw6HBTmzh2x9qqvaa0uNkityVRpxsHFBAS5kzxUwlqFLb+8PRqDTNHRXuGU23ovz4kQMpu
FBxDpw0Ha5n50LqNyl8e1VgdYuSyT91jYLFWE95W7a61+WG2F8eSKEsGQf76Qzotuy6lOcseZjNL
Ak+xbA7uje9iw7qsC5FBwRziaXi0eoJn/l4S1J2uXrzS/6oDP291Z7SLNk2w72wYfqHqPBXuA1eY
cJuK36FFbODGLkwKcbVNv9WxOXQnouViry0z60sWqA7uhmYf8hjOM6gqCkzA3G+GsSxn6FLGLCpJ
EGx/Al5+2uPxYrZ+0zDQl8yXJK94GgmTmcuakT5ZReHdaHXX1O3PPOqEAC7YZr7JdL3x77DS7hkS
N5R3bHuL4Vqrhtu+cjFJaMYXCIo4AatmLKck4Nz46JDegQ5AXZXmKdNsY/8Kw9KCocmnr36zXKLr
H1R+Y8rE+rn83iAwVGwzIQMkseXMblORbYELLnWx29ziSAgHn4XqMfdhZDvdHdz1ngZVNp9ZEeej
5Nm0br4isbUUtRJ2kk99inZ7adzAPbJ6HNC1VaH5LH7f1JGOC8nncgQ4N8T4qe4FmWHbKSD+ebtd
SeI3VsgZIWJrsHw8TRKdJJ1paH/65Ym1vVcYcvK+Kn9izDoCxwDpCqjSC86gAYWdJnqTxj1iJEjt
+Bip7EH/fH6sjjummBtRkrQnGJwTi9Uz0RZZQUBmmsJIEwr4sWKRfeb4damqpuEM546z12CxQIA0
JmaRHuFCoPil9VRsukV3ViOVRg/nL2Fpew2UBYYZWjDddHBNflOp2qcYFCC2sAiaCVrd3CrGjfLc
4hImwxqOXUdZpwp4C3HmLsBj3BT/ZD51we/nAiPM38EFH7E9Rb4B+N9j0Ktr3eRZOVEy1ffhvR7Z
xKhcQd1Lpf49Lbq3zWiXmiBP4S5GmHfyU5nVgJGxwGLVzqsp/gkTlM2Rws9RUgCcNyBHZxSDutQi
+m8LNZe1LCFx8kYY2wllR3oflDTdrLbnflW9XUJ1C30KdoM8JX1mqpevzevjRIqd+hYsLjGMTviu
6Klv3NqIwcPnDdBn+nUiC9gKQzgVmtjaoZP9oy+vOi5908dwKr6ifYBCoNOBZaFbWCFmdHlT/vv6
hmmUSGBk/GvYLKcCRme6bPAA+lV9uJW1YJGVdOpTO/laEUX51yAn0Ff1rVKZcRbu8+w48+nav2kj
4o4zJOCRxOuRhvmziPa713Cw5/Q11wrE0zj6aPJsmXtUuEkwfF4XtxiMguZBQKGzaeae7AR204Ho
vYMHp+Uyh6DbjzxE/DqeAVcggpmEMuKWjzS+zz9xoAi1t1cayefC6aCWcZupqT/arUQNZ1iwhxtQ
ijYSBbHcVWRXoJghrzo5FDmr1tP6JB4I5Rjpf85Oy6aB+HW6sEyyagg2AV4X/9MLBK+VAO4yxiL+
0lrLVNJPRNqcaBmA+jHtXRH/lF0xZJij2OUioFEeaAQNQKgf6oAHQ4MymVT5AA+Tf6C0i9agYKEH
0nF1uT2oJl3OEXEa7AT0ISyGlm44TsGHnNU+c/gl2i/6Co6YvnvRJKSlsoLZg2pudvcfPKnx7eIN
9jalfidQd0yd3FMRMX0h4SUtIko8I1uKMwKDbuoFkcScWPeL1AznWj4xeLf8RcFM0gKFpKRYoFdl
yS2E1HO+Do21cCagtPNL8HJfGJFoLHnXJleWM2MtAct8ycHXmWpT+0iJhNqw2LA6hgH9Y7MzKQqw
HW0mta3CagWbYVsrvjhBB+Z0I5PowXPF9h8N7LnBioRrlUlbyJ4sWHiev/VgD3lwSnpeitSuKFur
EqCaFjl/iMlYrh8ptD1cGQQp42N97eB80PsLSfYpSGz5nuKn0Zq5fA3vcZFjjgNud3eZB+R7R1N/
4pBxekk7Es8gJrAr0EeC8SI671O8JH+MhxTryiitnz6tBN6pUKVYfdx8fylMWlQRDM8awvxKGpLa
80qdCm2QCdBTkTg1/ivWJNZbLuxxXWT7S42Scky9utM5gmks9BaIeuATsgTL5O6THWCLwTotqCO2
QPC5yIy+t04K+nvVqcgxAM9i9c/Um9dPXvsaMHaYzk2RSCVq5n8Mv2EIn0+yo52NCy/Bsn/8+ilC
4slJfmzsFhAm2G0PV9nZC2PIHCU0g6flF9MG5hUM/Nz/n+1uNLrgcxwbvPY/EBYsM7NZZMa71NXj
jd9PEO5q69MsOCOytrPOV8tmUhkXdyE7AFtGCj9cNhQ5s2rY3qAWi2knNkC5Ci2wR4k1GL2J8yLK
dxraYNsdh/bBX4zndEy46x3Tr4HkUgRmGTvdPfBRZSublosqdMH3NWJeOAL3ul5cMe9ENNUacXGs
vhzTX9sJqabdkjjMHRgCUwF5rUhv6HRjBi4MdzLLpEITlUl/DqeYyWmsyBMHjWpIFTb5aL9irDHI
zZ2IjY8CKCYOrpesT6EANcnyaQeMzNotD+GLoVoai3QyXSWq2vxKmXjUhqv8VzvwBfNkEYf4LZ9W
5pa4D56y4g1U2LUVz4wXUr0vrXdSJgEcvhRh8t30KGd6nikx7ofQGlUOL/i/AJQ/Nd7yeZzRYotb
OSkWlGXg6YYQZuwWsjGAWepieqQdAA3GjBogPkwWDnAi3B49VJZ1jnf7g+/eMsKqCdVsHLIbetPH
bwFFmXyNQf6O9duB5stYt3MQXXjZGvOP9bVGzjd2+4fPedtGq9XMkKQtIqkpZ5rcq0650x5rgxcY
GufoYo5F7m/BYn11jtn0myCNCwZ2+OGA+k9v5kulUwfaJR2LU0LceMHDo+yqo1l8L5aHWNYhlqc1
6li9vSSiz+x1cOcISCfZN7E3X+LBDno3qq29uKbElt+sqhcj1Yo7zkLhTThzVYISJMaDFeFjWPmS
r7EngkSwqk9U1pVEZSM3N5wd4K/+uodR651Svy9Ku766dlSguILp7PA4XSelp8iXy8An4jsVI6sh
/WkunJ/Oe6niAxNEXYH6CnNhvc6nZsjMCMr97PVYVc6hDsy6wJQ7WEq4UC4mfajpvgqps8aDXF4r
s9/LhirhFl2TTJBFEZOtzx0nVw52DEkYsDXm3jYGsbKjonhVLYNyXU6jsoaC1hJHMHMJAD2T4Uh1
4kBxchJyUAcjGixOcyLMeN/mozEdmDfvC4SfQvBfLz9GuULfB/w608GfYSreb1FqgEcQCclR/Bf7
csXnMQLfCvLx0SFqEX1i+RmOiS8201UtXCh74AGoPZUbjfkaRoIyRJB/oOUjfMCz4tBRl/T+9zXD
3d4Adv3FoCgQYXjUXm07mMLFqKkmB5MhvOMty4hFPUiwJEyZJqojrdIaC1LAwoHiWp9QMN51kP2I
2omCg6/6ZVC40FdihLgJ73M0r90j3KhgyUsGhMLTWISeFQVsnxXyYWIU4zLbk4yF/eGjFbkAIrMj
IiDuywg2yQkYOJ1HT5/yHbzSqZ0AzUz3ZGoDysNuT0TT/cyNz0FgBGbXNkcJYHD7XU4dsriZMMDx
PdDTxiKTPfYEAQi5RGoEbZTEhOyKhQRMApoumDsvQxXU2fnZ1FtM4Hf0RzPBZi+5LvnqOLTuerDd
AsCu+J/ZT2enaXZ+Xr8PT/T6sit2VZokFnVzwTAbft9hBGtOEHv+bphVJkMu6ha77VaOuPuTPROq
zWFBQnZPOHfNj79sB2JNy6xEf8zfjf4d7LbSP1NBBUmrmAl3iRlxLoovhbbRjMNAu6VWdkn4xT0T
LNy2iYbUyxHbWMRqA47C+vuGCNwrALl2pHLtexdPcdvwN9p2msacANWFZ62Gm6vxQ7b+ji+skXGm
uUXJwxJQPwfhmKJr/CFiZolubg9LcJAkT4MauqJ29sDD8aauLZhaappFenv+QqWm1/8iYFTC0wKh
ELnmBZn5ve2JsPbNjzp3qL2UWY/vntk6oJzghcQ/cnoqQCrhm8IV92WCuOkrG9zX32qvq12z5Uqi
5ME8t0FSCJ95OS6jVbq47R5ydm1Gm30KoL7oOhtTBNS0Fr/cy+yknE073q4TcZXazBFZEgkfiU7F
i2NbzTqKGIiV0n0ndEPhl/xTSxhj4Moh2MSTnFmtmMeO8i42BKGju1FmjPO74mgTKroMgHh8SkOd
RH+ZtibMDx5TXe0utS8ARJpnN5oC02AACYo4J+EbJ/OL9un9ckQ2TpHM7jj7bbiYQJeXWu/fOQsm
t6rDQgf2om1PXpquY/rOM0ABolbYUTWcWQLdkbbiRPZxpqLRrf2SazTaMXQDSDsmtwwf8velBYLf
sJ/f26Chs3EISpMDno3HOlvLt58wdDq/biLGp1Em3/rOUNzmUjTX+tJzBijG03WZrI5h9IHMsUhW
3xYD8BQ8tcWN0Tness0XQ8NUbv3LyuX7YcNQsadDm92KN6ZSL0nqaSqm4ySav8FxgjoSTAP2rDhl
dh6NEmkh5FLu+B+xmgkPWHSlycPKFrjuGbVHDn+x/qNeC3xFLn+dNqc8ppB0xI7A4VBn5lTGlmn2
HhC9emKZ8L/W4Ofgiy6jii/poOIiKCuBiEdCIQWgJ5Rjg62hBk34FSQDhUF9gRx9WuzG98XW0Uu+
Llfiw7iBDWJrgZ4spnaOPHVJ+Y3j7HSGEJbzcuLoKTY4FB0kXErligStx4Sn0TZACi6KqXdfE6qS
LtVP5bEoURS27SHdhNbHJB8egM09AHa/KpRJShIyIjKek0ux/143A3EU3+PZsmzeRzMKo6FP1uYX
ZvY+1Ay+Wk1QF6xXF3VgxqCSV5j+BlGFntUTIPv3sWC4aMeAxllzVCEx2Mt95BrjNq2/0lWmXV5O
8ramMVXCo7ZNcFc5OAWpWpW+WoZEykHQ817WqAGDPxrrKwCDAEMSna4OqoyD6sIxOGSVXfPlnBP1
EfXQkzcVEMw2FJhMeIEwRxCwFYebiIbD8o2EWnpxWwGoHmpWmsd77/3u8ss6nw2GxF3pjO4Kh61j
HmfIOfd717azuXZYeWCXeQsSz6GsYB/3MIhBXeM9Lpcqs+z1+q7ey/YMfyPmchDkZwcJ+84VpWsd
QWYcoCN2aNtncG4fKBEGGoEJFBHYytPZ7PgtCC6Xqud6AaMnys3F8WtXJeppqGqMtlc04fHgTnh+
KD317/ezYnfX+HZseCOfq8Tt2MkAtOkdSGJgWoihB+SME4z4yUhQuInooihwMGxiqhxmIRgLGXi5
y0/aOum/O9Hass+yVKdrFmBsgxwbGSDUsVUn6jUsWESDYw6quSl/TkU3Cucp2kqmanoQPYsaB/0R
dqjUwgy79qhYXer2Uw7S2PUt9WdujFjRIc+ZnA0Fxo4s0JZ2W0V1Ll03h4mXfkEqWNDsL1JizXza
6KjsXubb1Q8eTXI4KkO+Imk5/BEd82VAIXoFHDR09FBLUyEd4MbpFf0ASKH8SJ6ZubTxQ50WYCGO
LqM/U9w8VT9fNYe8lBUIKU59BGbqxkSY5eWxKKxuImambVtAE6Sbh8lcBIWa95DT31SMhD5j8NFX
nLWweigU+kuIahRKSFgrdDO9mQu8by1GdQeGAth3qSJsS2rVftYeKjeSLyj1iuYNHuDB/4JL8W4p
HnXJyuH6yzbldG9NYTjJDvwSjkUm4/yskcz7APesJcbkfXsa1aaM2MMMcJjvuvQ7MAJ5KsXYevd+
tFqTSCz8kJPNnOB/amAw/S6X0/xEaAeR/jH0wSxx2qoyAqIJcwfqWPDPOfMydFRUvv+SztXvCVSD
QjsoGjKYV5BrQ+f5x10G4kxV2Qb0ls0uTnSQTZIisYqtK04nP2AgC68cjDmqNhR+MKNNwJATXkOB
FrmOcwLyg+/8i+dQHFgd/hn/ZiBPUVI8lH+uhP0A6w5TSDgxkPan7JqyOKhxGgzHVZJJL0Yl3xHR
+/exxjZPnblguhL+nYIk4YAsFn1QsY8nDjmxJOt8ahBkRB6B5vNqK/N4crVcwVMBLLuZFVGIkyJV
BOHj3vSo5ifvzRVo3/tKOHiwkCHvskOYEjdBMcPj9bre5llKcgsP1HCnjT8yoBBIR5oAEQhBYtJc
r3W0+rCu+uhW1PMC/x0QsqHjL9C9SEXASIIZJgf0Luan8xVkZWKLdydzPfN0mPu/REVHBtp4MhiM
wMfIkE+qMXsslAt8LgZmS7qDJlphh4mplRoLJcCN9vdJam5oxDRQprNbRWyKNYJfd7btZuOrOQTM
SEkMGP8zAI9xSzaUP5qtT2S7FGaxD4SHaPf654ZKVfwwHzsCq3f09zraYH2D2b6l8/s2hXQZI9Rk
zjijvB/gUn8kPjzqgb1dqxl9lzIU3a3XNjqpoRzaehMlBNH9oi+DcRIXYi9g9DWjL9HlGKgKkvq/
iV/mC+AG0P6wndUStgmLJGi/R5Xdm/NAtTOqyNzXc6P+qXpRiMNXxD1pzY8Qghn8jZoQYpr29eB/
BJA/rulUFbk11q+1Ane51zUegS9UAb0QEHYGHfABBXMvT86EUC/MHMTbWbcUsrkpKFEXV32KAaPe
7uwRLXMng3IOgH5G1xmqtyxiN2EdZd1vE4Rwa1rLl+mo7pxSksdpWb8vBmWfG5H2HayvJV7EbOkQ
pGg85BPiqqIaGr5QGj3mqvSIWC5Yx0QYlCBB8WcSbrX9YuAYInswpkbTi+OdXuV/0MgTCO0t1G9n
FbGzr9katuFtYgU9tgtGie7SMpyiCkisHwYb7ZUXQXvejemn+gcp3qN8rETEGTz9KPlK2hZi0y+x
8oxPMx77vnutJ1cVT7xcQIbFTnkp5mve3en1GBYs76FOPvNyCN1n6lmt2hsttcUAqzRLO6p7ktew
zYCukF4Dwmts8AI7SFLcJM+eEixCWkRqfBwVMoY+rNcAa97EPDgPU3S9n+NFVMX4cqzJUwqrYFqF
u0OuIkeBUGa10UgOTYzFoo+YhyLUBLNDjmpej3jHsfgqjfqm7v7p0rchsrKxHLHEoYL4glozyjvE
nps/zmV2uUeL5056n43gTmZM1GO/Gjkrt8wLl7ihvUqvZ8BsKIHqQ/20VzfE38kZyvpFVqBcf+tQ
seACRvPyj/I9CzhwhkiqA9RDe6gw2nKIWmzPYvPkeVc9moOcObWObZfUpZSb3kbOplYX/fACClCT
yWQVpXyZbtILEf0wSKtO0NT8sUtjj5TDxUjb4B4tpyRrjeVtbtncN0StEyRtzFZyccA3UBe6jQgm
xQq1m6iduaYPPPqErOo8j4ew+pn5StmiWw7msjPkp9fBkUXjXVUMPoZFk1l85DhRHy1ONw5D7lM7
7vEExgzAJFKhqbOVyLBSaD39N4W+EWSBB+Da4qLA9VApr4+kb3fIWh+Qvw1d8tQlygbO8hAtB77u
t+t/QOfL0qVS2iz5XDf/dq6m6yDcZacUeFaXhWkeNkbEeyPC1dmH5ZJGOb/3wd6RJODGFgc5Td55
yGphZjfNOjP0DwBu9xikSRBGSfW2nkynXz+KkU52TgR4G9zDbdE7OCIUxNuO3QURYr/Xg48X3sSK
8wFxHqJHvPk22uwULCUjfrxclA8O1kqyNBkSKxjVFuHo7IEFncGTDO/xYfMvi0THlkxBDTkhy2Sm
UJeBIRY7mmAYCrQ4woyDRvMeirAJJ+ksIxB4DWBpBi9RyXOUHfJtCkxtfa4tMdc+9DAvrL+DCsQJ
eTFeTdfNw3Hl12DcOBVuquO7xwWDsGGhpdLzO60TfVdjZJHGUFkI1FtY+FicvoukVznzIvGuq6d8
p9FLru8mk543EGACySfp+dWbOyaPabfM3F3w+Q0Ua1gCbxsWeYBjCmoMaZOkgQqV1rlN7xdNLuhW
01xBYZ/e0udb++dmempHAdXMdaW1T1iScWKlT4QPzKsVIFd6ZqatXqr6MirSd9IpQzMWDC7JGnHY
KDmsn4vJHBxb3VcDSWIUK6e7k3qEARpjZ3h3LnE0Ju86Nwy4eHHkEsC2DTv/YgrtZLXQzdlNCqRV
RRBP1c3+ZfIUICq4KtCbbPtTFGYbWbtpbNu9ZNX29LIw0VvtX9PotvirmOnVdyAez4BfuM1cFEXR
NRlLFaWxSa0b66BBHFzPVxjJKjPzyX4yYkDEmvpE4ikPvgSUYUtR1OT3MCdKk2oEnA0yidfXnZEa
rb56EA7iChv4CESLdmmV4/BoAkXNqTZ1iUBjyfbhwfVfDSEJJOZKECdS7aJfd31O7dRrt3au+uVs
RSn9DAIEJvkG164xgy5nIqo/2BZsNMOds1SAcuAti98itPzlAtJ04VMKm5uaH/vYt2MNVvEZwJzt
3tPsnb9Y4iuPCAYSN9o1D3npYqdgDeVq8nVDw5JiuS/AEZSHEaQ09erEHabGt7xyv8qX35muCh6I
vfINTYR/a+i1+Zjo5kNfDIZYipYDauOAIaNlk1AZWL08+gJRUMh1OOsAkRHNTN+L4cpyjb1yra2o
BgY5J1gcbFW4vzSEpERZ489o7pXKbAet+Se9ytNlzIXy58wSDfu9h7v3RyiuB36iug5SVNSPs6qT
L5XjBdWGz4y5opmExRpUzbJ7vyuSPC+Z5f+PFvtTSuAgpkXUtCsto4oGCl8ImjkdqbxKw8aUWzkV
zoo9u0Fw8xVmVJN6b3+0hsmovv5KqtTNMDrfmuifD3X2/S/9ncSvKRTahxkiTd0lWOD45hU9WKmM
XA5F2PYjk71Tn+72j8bx2EhXMx3AQk9U12ltCK0qLzDG+KJiub//f1jsH7mo59rDBsK4YNsSUPxh
qUNSA8kNJoZpDQXakzJSuPo/4HkXY3/w9fLgGls+rHS5LGzLFnOEH7K2JNzCfaLf05E9Fo1slWEL
PvxLiUCbbwtP9OQ6sAlvb1v4WCDgbIAXZtz0o4oZQ3Wdei+ZIGmpdZzEGz0aUhA4JsnjSEIAZ4YX
jZa6S51d/snZYfMdg9eipHmjlLcwrJTiH9p5ayB0pXn9l9rqEEqg7bmFqi1SFqHE0M8NmoHzL2Q+
MLJ2UUF26XQ+Aa5dDvRikMefavCNjoW52yYcJLgQQEjWJvMwxW8ZWNGjoPhAlIBp3C87Ss46MvD5
LWC+cEthmkBXKtPvl/hxEJ3kqIr1YKxyZ+N+BjATFjAjftX/PL+zoXGn9t+nK9vaaOfXkKpO2yaC
DLjw2YnWcHA6sxL1Evi2bjjlYix+mXqAAMc4r80bRmFHEu9wqvYeCJnFzP7kWoAFTudn8xxvcpDv
6ocHFi5T0ewRn6DPe4NUYuLt/JRq5BBq0nFlf9legTU5v5LgC9yrZiQ/QB7aeokkpOYKX3GIxxKp
+Ru3BngFTqWnrHipp4PV2XMw/m8XEFSQnfSDmHLWqiHarLkFd4r+ZFrpjywGMEKvnS/uJRJSvvPG
rHeC/ACNC3YkDylMU7U/LjindY2xuL1fWAUIC5uJJ0kq8qQpb6JXT+3vZkziK9eBBIxxyZgU/Xh3
ndC+AxuM9FTUxgVXpqW/jb83cdljCRkmoVvWgl8J3LV4ftZiYKfWuvm1652ASR16nZeciTQVAvHu
CwsMVYSqv4ExTM/lgLPlYZQrNz0TH0yn/eMGswq2/gdK7IU61tz3YPLMwZ185Ve/PgpsId4FGyQZ
MKhISwPH6lk5t72xEyqTxbgD6HvXQWcSXqjBc5h+s//zW3LAbo8hd+GJF1VaUqnLd9NZmIGU3BwH
TauzFVhztw4BHmiDlyDfjJO/Wi/3IuqxGg6OxJ9bAVB+kkgRoqB8lCr0Yzc2YAsv7jnSPh/THmuQ
F2SNogmeDW2cEV/nkk8h9r1irAG+kfKvEk1jLajT4x7pzoe8AbHzKdmmnWmR4RWBJEqqzdU3Vemq
6MpNUYAlecoba1oninpYe2LSyXvLr/PAGiCKR1EFOA4/Vd1vMzhh2Z7IMbQSqjWm/pATo+ChH4ru
IagtJwAi1HmUwLZBrlXvxSEHPjdYfdPXTUEbe0FXmuuxJnbdKCZQqbA+bXzriF21pM5x5BNTILio
CYGmB94fZPoTGSksy1qzvSoOEVcof2YkTcFV/0fkgYv6vp+P4n9bM4BwIVpzEbYykc5tZHp9i6tu
EMnjI/bsE187Xq9K0f5aIIrCUQRrLKv8U19dD2uv1UKw0D4MB/slLRppyBXYCe/tBExYzOxkZUmp
T4ZlGNpPlL0ExvW0tiDylAS06SN5Ti28cvXZuecnU2zLtqmnkxzAAeXkHYHxvc20ZvWK5mcOR4By
hYTE+s3/jPd2/nT04p33DR9rUUGx27blYrBBGtoWlzhr5JQ/ucsFiUVS+Tspjfg2AZVJEOxq2UpH
1gln0P3l/P+B0671kkPAYJwDKBoTBMTNE3WsrPKl7vgT1x7VJvJ68TW1X/INMFJJTZyTvKceOsMm
cNm5lqKQdM/ex3b7HqXoG9ASZUOtS/FglVkHf1PUk4nxplXPgy4b5fPQv6WyxnItms3hovA302RM
9SAajnXSac0xF901zCpKBIfaW3zwvcFggIvUUnKIcfbJUVNcvxnACheIb6pLClLTs2VcqLivZj58
DCLzFR0PydVJTNMOe5CHWpfqyPU8P7AgR4dED2q17L1POaG/NR4xz+ddqMvTcdlEG5SsRiSU38rB
xptjkG4WOSNXja1+QG3T4s3VDRrLugEnLtm7F6t1iErxgxxIuqQHVE7ehRhV6DXzmJ1qTI4BU5/g
ccnm3sYUqdfW9REk3x1nGC/cxNKIOrkv4s7aGIMtrGXc4rLkX/w7Us5qKV6Kncgn2OA+PNOtTCYk
FYvTehOj169x7/B8GkKGw9u7KwmrnPL4LuPmrPbKQU3lJJDKLhpG0iTfWgJUyuCBD1aK6tuveEQg
4lM2V3MhzeupBysmZSavYeuz6w5WMjqESko522J668GoKCTTTYVsZVWCem15azjs2f0GoqFEwzI5
jY5ak1J8g5KnGZ/om99TQcImN0+zHRy5gb1nqNeK6mgE6M1topwtPUpqMjz3nI+aN9EDzNX34OHC
KJRJ2U7+OtRW/+aj7oBAsxjmEpK11zcvBHbl37w7nEfZJ/chh/YpwciwPXVkhzbuutZN6wxnVphP
IcqAvypfYqua9yAAzMT4rL8z2RrrKyxngZoZ3yyMsrxwAyQ5joGldY/CnA6kD6T40HZl6YdxXvVU
2jLJWErxDe+b4pWHj+aRp0JN0gyeyxi4mzRNG02+wodwOU79bCJ13z/MUwpw2sDghynvSqRSojjv
0+B4mPT7PsvyrP7C7D2k9/x8v0tuxpDifXYDsFkJ2Egb26WOx28iqCYju68V3L3Gaj6WUIHAYzIs
pN/NNwEaeOXMjvUJYgXbV6Mu2QZasmW9hLhRpnZTkJYrtABMI5aub6CdWGnMV9ZgpsMk0BDJfal9
GdvWpGIQXyGCQrQZZi/cDgnaGFf1N9hoQ57hTkvezdDh5O5J6k+wU4/UGV6YBYOun+6n1KOegABb
ayCE5jXVlV/pNjoOFeyEM8pufp1gbANUgUmo7tE0KsUXuz05TrUgtjQ4A3AlZAOicVPvBa5edWcz
m7O9LGNW8HJUU5FnGOI09GPjLpNDGRfjvPUW1FtWQcay5oXrDcDcAOw7Xo8iAzgtRJvbSgOUtXDo
0Mp/7kKKryUZ3J7Grfa4oqTQNpYMqDl/yVJVFGAq70CIr84FCROjVsXBgsCaHaEuccRV9M9RJbmz
rWHAC8KD9dB1UElINU0rHfrgi/qQKjZcMT1FtkTsfXvKLJ8MdnX5jx23snDmlcmkvpoDYlvyGRWf
c8PyLSKkg50IukpE4ORygHoambbRDTvcnCuPt3YW4eOxHxpDW9F+lBMkw7Bys4dD6XcYcJN+2G0b
pFLF4zUiVoez0ZLttZdR1cBWAaojdimrCtnp+t5H8PHcI2XbVCl0JV6mRGq5lCs0xKpGrSEexweG
Qfmkd0ZIqJhjhp/7YVTkkEVnny6FHmSr815wg5bKq/J+BDjLtmN6s8wNEaQ8cs4fzgQV8HXMkvKX
y+L/7OxiM2HohUSkiVCacHG7nb2UXUgYq01TCvfozHHCJbZ1yPynRfyxVwYhmU8lae9VJ/DLG0HB
ehjdd+VkTZtX32LRvo4yWyustN18qZIhtrMT0/WDgAUBCy5N99j5lJ27xuG+0mBDEeaIsGDWLBz3
ZCgKAUxDMUaj+CoWLXPuVI3KXhKlx/kcjbRyzIxoe6SKXcknjeNG7chntqR5Xdf68ABen+mMCphf
xJQWVTE7Ll4l0LdXkYA8cHFEH1WA2fXdrQ67uCyATJTAlX470DCWLSpmOvgN52RIMiAxxZy7B0yC
C6Bb8BDUN41rmMQqTs9EPMhmILeCa3lnbOp6ho7QQW+SKDike84EhGJYijFMFxcEvknDQb0hunHP
Jel1Ohj2SbMjBODRshZeJ2qTuobsVNOvKWiNr8FyNAxm2BdqZWKM/QTNiM5i2KrDe4/nulFo9PoZ
jv7Ew0a9xxMDVpoSO6vkZkKtKKArooEsvG06b8ovG0eIFt93TbDnLxR3aZhi9uJ8W/194RjOZ9+y
EZAq0mT5rqUCfZTVnnMAMPwCia/hF+8ga/12yvZk+EEdOt0U+YXGFYs8TyKa8qN/aNmG7WEz0gP6
OL1i5uOz2Iz0fFUk+j1QM9qS805Uw4sFHnyDoxDhkBPkcfIhOyGZeO9wxEcQE8WWi7vrIOfmJVbd
xZFzXgzSrasvMnt1rw2anAem1zpqcgcc3zbqwzIQeAJQGX0BZ3tSrQ/fLQtvseDmBRNbDTvJfult
AQFJIzXxXiAgAChILjx9iaEe+dzHUsc3nNjPe4y0/FU+AtHt9xyCaFRNBMGmb5wlYuRf2hhhJBpy
wJnoNPpdVocQXcD5OgNZBIzzHGVb10qZxz2KDi2N78lBOSM8zD45kFWYaIGUA5ro1GuOcBcClp2r
lHw2c/FkXY9fNtLycU2Iaj4Hw2HXsd0Tqn1pDbpD8dqJGTrXz5r40HVtaJIftYv4TrhEO5z/JFQx
+3+wAUzoknC8Y+If9Q9tmjRkSDcYKVpzEsmD2KDMpwxvezH3QYzMEMK2YnxeJxZiRIWvhPde7Agx
RKumzdTFlKUehk/ClW9HmL47324iVB9j/TkrCZvaQj2n3G0vsikMEWAvQiiFItBy8x3bLPXVp8Bg
TsNDfSurlyrBMn+3IT14aWEmc7n6+XFSUo/JiZj8+FXSTWJH8KahzcpSm/+683DOPQtOb1UGlXE8
WY33ckQJ/MRJLKt/68JPw+hjPX7i1OkOAjcSDFg3dUckeZiKWvf8rJuL8347P9fhQM+jkA2+ehEF
XQv2bOYW9A4fTyOnV6vFR1r7cxmM+nsUtmoBDApRMGGRB57tLHHn3eOCCdUuigDHi2juBwvNeSGn
r+pc78+ypJMno2pcZBQnhcIwn4tqF21TeDbaPgRpc0uzygUbtHjeoIV2aYxDBW3zw6nrLaEjizoZ
f+XzvzYb/42R3abIz2PCWEXezVDiVyKV2qXR4wMFZ/K5Z1LyPpn5sn4/qK3lNOpysdHqwIhEHM/z
BOgpN3NEJAhegKhpdy5eL6hMJL908vFYSvicP/SfQ1A175mL3AL/HBkgoc01Y4DJiK4lVfl73gh/
NOkh7zmuMeDUBRd0gFCteYNCL3Apm2X50okHrFlJ9ys0SLPOyv35xWX4ILUeQX8+nm9T6YFGSyp+
p0pyevAaPaTqLpR3eAkDy2B9jJTn4bH9uqINtPesJrnrjeS9lNWaxUSE1ivcyX6fPgRqXSMsEO+C
PAwB1m5r8P7SNUMnz/gUb+iU1qcRliC0A+S2b3wJAYTthgsxuTp3LDIZdW8IElH8GqrUBcpbBGZ6
EyvCdkHiW0LRNkFikKPONryRkLmrpVEwm9oJFk9pJNxQXmhvjVgVg8993C5QCJ7BPmIj4cQmiOC7
2j7xJ4Skweh11zAsVt6jIKk/0ic2YHJnH/ax1rmY757hOXgkbYdqMVyDkbb6geqQB2vTxdQ/RhEc
4TjcpsLyruH2FFospIPRop16TfiYH/n1kd0JEyYCAx2PdOyLLy6zKcr2xz+GCe5jSdViJyRi3wA3
p1cbykHZ1NUy/xAEZNyf20DUuzbCAX9SlafJOVi6h/2edy6qEckV5669lGWThEH+sktmDKd9FBR9
mtTVp914M0UIDvecZZl6VrdY/WhwTqtymIUG7TgCyY1pdgv1AN59Nar5RNuaeUJ5/lsPspK2Mpe6
y7KUzoHKDbG34YqXGtld3FeZAAYkRw/7NnEUMjp9wUiHmhEpeqfOFo6oSSv709KudnyJFCFlhaOd
FJmVQcOx+7SJ4ZvgHimExn56QfiY1OlUE0xpD5MbfQtc3gIg7yQQmqXuCMZz28b4FREnoztuDDbr
WeH8+YXsM5DKRJiicZwSaTFnxSr0Httu+/0zuNRxykYlnViDqW9ZGc7pzZfWAIsZlVbVlO61sW/i
aR9NbF/sz2qm4BJc/mQ2ccek5ztgQjxglAfrdAccNz/lCr1A6+K42Fi0oiOUVE0wwnbl3ZXtfT8t
tHwOisArPacOQwT7/txmC4+45ETPQEdbltEhZKGByHsy/gkP0sDTd8AIOMzpjegeVbSddQEvUpBT
ZjOQU3bYysI0Ez+hWga8ois89V87YVZSQthgkf2vPTo2X57Mf+igDTi6DfoNe+4w97Sd26g6tru4
3vlDyH0IWg4QW2TW2m5ZyUq5wpqWxobYhyJd2dP9mszZjB+Fc+5+dU1/Fo2a6p6390r7dbV5ddNI
M9Io7bAn+7fM5Ok11KJ1yevbpNzO1Mv7EvwolMRpLNP1pih4tU26OvdsTQlvydwS/DypDjmDM60F
Tm2nDxNtBewzFrMqORcAHBSj1+QdFAtkBrkU0uhavTBYi0yhv1MHGAvfE7SvQBh1gz0VebAD44QM
YxppIzDV29qZzOlJ0nx6vgrq814CVc3swv1fCMAs8x5qBKfqOtGlLKLBG7cmlDomuLyT1RDyXLhl
a4VJIDGfyH9xh72zzxZKTqy6GijSM2bhnei/fZ6uXgVzASvxOOFM+KVLcsycnaA8EKH7QiS+mZ3X
qy30C1ZMSq0uBUDO39iDYtiH7OV89k5iaAi5GeClAbPgWvVjReUV/FhWpgRwfWcNgU+jAFc0YNDz
/bRspdODUmAi2RGja4ILKLDVCEI0L3y5yGNJvkfHXhPoKF9650lwTL5JyjZKozgFrC8lKT84hq1q
ELtgcj95IJdP0pqoduszC6Gu9Ivozw15GGBBn/pXfCatPqqpjDuj7O7ZCRqBUQRrfPF40jycempt
iophZCr+3N/Zg20RWjsbd3vbANJs2wY0ivNIFNzkUYRlW37Km3YMDJ0g3a/1SwFH8HWVm/Wva0Mq
XFkkGQwHQ9bdUnLMOvxireT+bBWut7O/6Dp9Rbfb2I8T7wa5mKkP/erCGgXUXWvA2uhJ7GS27/2g
fAbIKGqLZIHvtme4469mDETtriHI4eutk7+lQ+ntIHBMBQMP6nvOKD2O/aVvOaP6+eLPc4GxD3UK
gFrH7dBGn3+IxurRyW8nBQyiKEvICXy95nkNe8f/QVkwIynjvaR70OS04UeDhX6e+H/PXgoJNDRk
5u/S6jMMpr8TswwXVl4Az1d/04EGxEtcJHEjBXWFNCiPXmyAxAaEzmMrNpQsVdpEEs+E8jQpfmzZ
FnU5r5ExQnKxpARijmGthCHalsGPL1v6v1uEvT5wp5DrHlWkonje1LudCmt/dVHNriGUCZPUoiEL
cACOG1KqSxfXrK0pnfPogj2Wx0opXCQKCAhao9EqhsmbRA3DnFGr819krzDeUHG0nw3gQiSJPbTM
lhJOjX+UM3n2M6IdaJtCl2mQ9dzC94xv1tqfjJLFMZM+l/ZAgOadmPJB2OsKlpKDiYjYSwGoGb6b
TR32Brcy6lbw1o9REwXj0740qz6Nwa/5O386xmvtleQGCPBnUCXbGM9qCV85gXqqxzxRPP1pMbCe
AvNrbxBUM/B8RgEtzm4X6jwE2GqY+3VtwPuiFDAXwWuWPlMfJCBOD/7xiN1IQojBGAxJfu+k/0mU
H0VjFBtwlfDV/Qze3x1sJ51eSsyGuEcT1jLdtqGa31aMsItgWOEVpqCiM7hewfQz4gSP+vXSAA3x
X7+xu9LW3TAF2DQ/ZhlNyVZcU2sai17r/IHPQH3GPVEfa6X0HRkA6lfAie9vEScrM6Y9J465ZO0K
VopcRDog6SVfHHmevjq3dp/PG+Z2r4qyOVXGERZjpih6xLYpznkUUzxa9zvrSTJmWV/8O74prlgf
7P9OqgK8AXB1kdZIvJySgbWQyiuMlYy+Up9vAc5C2g3qDSGJwT+p/RyxxDYhKJUEN8HgI11fY/EQ
LJ8NdEypzanrCUiFljCeD+9Vdvm1GonZsKOpUEgmsfpT9VznHVLWN66Zt0Lw/lWGaKxsDU5x4m/3
GEk92XzhQJJKU6XuVfLTRXrP7I8VX2XIeQoUVWz3ESVB3CS9GCuuF4lwQ7GymLISpaLWob2jG7H0
mwSNFZkDKAkdcYe9p3BpkpWjpin8Bf/IpUhjEUCoFbgjdjCU7svJxozUJQ9nK1MQ7XMQs+SJHBi5
edAvbwQDxLB8j+dJ3BWwIqycWNErmR77kHHmdQMzCIRXOO+A/PQNeX6qHHfJdz3LKQKUykBbL1WC
x6cGWnZv5W65GjR67SthpZUMx2zqe7ZywLzT97gs91wbESvVS/9peEiaTdkW5Dt60OQIyDqt+jA7
myEnoQs50S+ia6S4qMIZy6YZeq7NfgGuk7QzJa+jwSnS8m4joB0csx0tejtCepn2EewG6t4XP/6k
cEHcPiOJ+YcI3xn12pFJRJiRloHcstsre0vAXprbVJxny1rJshcz7l3OP91RQtzcceQI1TX6McEZ
prkgc3pz3S65XA3anHU6DbpU+HkjfAHjeno1WbuX9WfInfrDpa/dbkMSwGMCiAYg3j49P5BI8/lq
Qbif5S0YZy3wNooYDC+zsz4N5tDO43BCGmhdW9+xz+sqpP9XeY4l1VfxJhQJGwygzVJb0ws+3dV8
o5WnemjyqK1sfHdBJ7VKuHMYZCaN5LPEMxDDhr35v2IHb6ggV6XQbaWEtzWZx6ZNcOa1xv4+vfv6
tF0PjZHOOw0ysHFydcYBjjvutivRQDiQIjv6I5d3u24SLt0CQfINr7RjabIWg20sMShm/a9ouewr
DY9OtThiKX3qeNcOjx3sTNwrb2aoKwecKEF5oCRKVWiHKeezRDlZ3JmoZjW3+WqHihxAE0pz0BIJ
bfoCvUpXjYH3cFBr9qpjzHoanQ0YKYluAZ3N/z5uxssmx0t9KOp4YY8Q7oJEwH8mKgerncZPUdeh
w3oyUAtcK7jPkZYmnQWueKSlCCaDfSpW9RTuuDe4mskfIpV5ZoUo4DK1RmNiVb8xpzCxNYV6HwLA
fVdgJdQUvqJHdw9PZF7fvxcDFfMnHVjCpoGzrOOxyWZZPTK5O7El3MyLB7tVKIPG7ArMngVHLl0o
SSXmWNUopqkm3jUVsYaRd8bnudayugYQezPI5b0l4tREXFf2iKqnvGYJN770aqEheJmkHUVedsc0
jt4PJhRyd7RwmKbI77QRxvkePO/UUnN7Y4TK04KUYCTJgxRdOsmX6w37SyFZ4XnRCeihIv5yyfeX
88ffNLhuqcaHrvDEKQ+qZ0lM+jbmEfjBqCZlzRsWjtOD+D9ewBQ62POitrJVK0RtGe9+pp9ERRDU
OELgYWoSWiThKVDM4M7jnu7CHkQXG4/AQshlqi+52nXLRxxDuacqHYg8MxSrx0pDajpNkkQDGSlF
ClerqoSIvSezG9fEOgfPWaJXrpzh5BjqvRBtXwm8bLdjMr+fxlYgHHay9Ut96JMfHHzHbhgs+l1C
gFBQDhY40eebf2TcNAHa4qFeAhLonBDowBIoeBH4I7tUW7SegKMFPlLEfv1G7rgHsBAI5oyaY5gB
sGeYq6KQWjZFv/dulpUt/SB2m6WlkjeLZFXrCTOZ5kxTGpRxTlAT9Fe4OIN6YXIYPRkwpJWqQChK
AXVAPxxDdi3nFum8IJFyFx1oyCpj2lgoM/fYx6Y/lR+tknvQ5D+6olhIV3xRR/j9CxdbgUl7XlGW
4ROmrog9o5dAOjlVAj2WxKyUJOocA5aGwSzOLvQW6JVmYucl6TvYLyLOReNWae1e40UGVPc4yL22
ReivUMAG23kNpem78ooWGfJj6U4/7bIwtw4RL6MfNugwbD87s5F5cWduU4/LeD6H+rSlRzcxU4rk
TdiPR8U81u+vMWJm72oZLPRa0H1HjVvIQXXArxmX0IhwtvkkT26qwb1wPB/UnofI0HqNFP77M8td
Uepu00YQ19ufLU3bxwZRDF6Qn6QRcapgLgbMKI31B/0pjT6X7CdU0JbxpqfxahJi65r0WR+Sf4tO
cKVjX3Bnrt7+e3OM6w77Up7iQnIN2O1AmJtPP4FXM2ejo+b27nIrIsiBFvawshQXC49eh30JdrbB
eKHklzk9a+Xfv7t30iRS2qkzMiZQ3vxtqZF8KhLCQJpOjo2LzyfbYc26S21Rucy5E47D8+cG7OZT
FKA8pCS/N0jHuV7ECQLglDl3UqSta7jxdAdq5qaElYdhvIvwZ5mKAtQOUebryVDKXM7a2lwfmmtp
1zZxXTFo+7G+caIvO5PfJh/skrsJxJU/c1+YYFb6hRMzJgEtUxPb8NwG9LSYmnsDS0MQ78bgYTiS
JkG4fDj6/nGoT+/jf4tpyqvHGlQakd8oO6/jZtqk3uCjwEbyYoH1nluDoGPq+r7877LS4yG2zrOc
dFZOTLENs1Gu8ZM8zmvFSeoUAoxq+NfqixRWVadEllA84JwRYlp9yPnQOyc19btmo3FqDL80rjnj
MoQ7paM1UjE1JIcA2P00od1lNyxYRPfzJ4J1bIKucE2DyH1x5mFkj01n+rdlv3rlUYMEDeYTyTS/
APjz7ouhV8lpecPBMvB08XJW5j7OBIosE/0VZMeJxGX9C3Zcq01rcyYCxo3gfbc826npbJtNl5n2
lUlh1q7/kOTAXuJnjco704w18QOQA0tOgjWYODMzSVLRYtuX6bC7ulP9F8y0bjwwPLkK1MxLLXz4
UNtGGEycPDjKpiIPGu9oLMPRX40iVTe+8fE7D3yUgjrdjg1MTqKhYoXoaHYmSQ4doL56U64fWw3s
6A9ja/Tj7gK25Z6LLkWaGYHiGg9/wem02pp3C70yvfNr5it+BtCaNED3pz8SSqqu0mP4sK0Wl84P
ZvftmuxtNEYNBWKrEiujbIWtcsq4lb/tnxKlsOoOb8RjHxRNBRcZiHarUuQS7Wlt2c3fc8W1L13/
Df/fngQq7QsIN2AI5iQ71u1H9gPU/mFwUmGSPgAN+i33I7r1QPm8Piv73qYqcs2+R3Tsd9z6gExX
USzVyd3NbtdjA45G/ZezQCpG+Cljj5NxOLs4HgrnHsemu1VWbio6F4CkibHsuVzdd/RUDbbwpjpL
k3h8AswzsYY8uMtD6URYZvNGWPNwoQJ0Ymvz2XFU0AO2S3w6FtdrJWY7uOYd4lZyZqNHY1GmygGW
GOawGBhGGHlh987aaLBzxfv2a9eQtJI0fRQjPQTRQLboDtV/6lMLbK+Lycv9bhsn3ieCEMdqunEF
ceernZgiLh4b0kw7E2HuKOoT2EDS6xTqc5fPzL0mcz52fFmUS6NzMQ8FAZ5quli2GjtsXH+Hsyhs
7/NXRhZhRctzlhrW3Wj/5J2K5S7qWX734PdPlIXxR3nzeg9ZbyD7+qUTKyrqACyFQ/GyJl/zgZVX
7T365HzeG2j6Br3cMydYrxTXmdwgwouVGxQJj+RpG64eNs6V0Xb4rhPqdVV7Mq0iUlBufrz1yC+o
30/UP2P6pLGTMIK++bdiCMPYZYfrcgiDTcJikps3v0kwN3I9DwA3CnM0cy6HkB+eOauP/re4r1qT
SE7Cv01/2QBLdmG649xZO0JtyejBWfLU5GW797vCJxw4ul2IH4205VtAqEeSPRIEmzVY5i33aFkL
IYvxQD3/nMmxTply7ItAyilOQ0B4yN5g2I1KWPaX6dPkqIAYKbYD2h+ConsMRHO6fE4RN2IeQpjM
vZnjlfiABkG/s2OIRM/sTS7muZj+b+btR+mDhtQyNxpplFwUsiTaoraJIHUwVrSBZGZeWLlx8V88
bi9erYZsQ2D1KbLt0seNq5pU/naIjt5E/wLWKiRPvKTrhf7+utbNwzqvAbrjROZ58GV4YeH/WnqF
BFNcGtW5K4ZrIXbBYud70Ih72Ozn+WiHc1VwJIVHLXmZoPDMcCeff91/VCv7qzebzPWAcLWne3eL
tYM13p3qXK5jPTTKUIu1N2wyYnpRUxelJXnY5EgNieUse9e4+ZrJMCQ4AM2XurhDaAzK/HK66GxM
+kAxK57YsgOlfAlqsgbw7l/wvSNZ3BEOa/f2aaYEGM08FnwwvZ0EQlzWffemhM4WPCJdkpFhI/TM
yOxYB6EMof/n5d8SWfIki6bzxMmVleRIsWIsrMmPPh3WepSd6HW9q8YGHhOYavnSrqk7wi46PeUG
eg32TPHknU8Cwdm9PC4dxpSTYCY54u7ZTjeQm+ubFFS2lRGknmVfJCae976aihj6lXpaYh3fUNc7
zIQqosi4oYzXuJoE4FztMaXDUZJRCZqEednCzGECstAT8L/Uz6G1POLBNcEHaCaUlXGuraF23/jF
v/au5Vrhi5HUbHcqplOYi6ZZLfyCjSONfPXcAJjxQIt54oxfaN6RSCIX/ODXRX2ysjLgjDRAhQN0
BAO8ZAZ0gYEtzYthXSG+sJfWW3UvWaObMQHTcTdykjl2CYig5G2OWfXqwV/MsXn4fbLoWJfQD0XB
XBdCcd1OMA3hZ0HA2MbS5o0xxOZnpgpvawjBUjPybUBxKXVOUUOnAcVitaVs+TZCO1gxD3Be9Vl/
OUx+61Hg5azNaCGaZGxyM+tlpo27nNp9Ec668omQnWUo2edA4QfoKJR3J31FvSqR/dBZIBko1r2U
6WrO20RaCXlASpVNPCkJ3wPmQE6QGg+AapHOLXSoZRq5+dyA4bV641si4z7qvdQU+vNzpCttMpAG
7o0BjGwNf5yF2VjRo/Tq039hFldvu4uUXEGeiPWSAbUos7wvVtbHA7KnKFNRMx3+OpmgKYP0gCvN
ysgRabroqfVs+vYy7xBnRSm0Vmn9VpgRzW7sldZFSbtTk8TDJDUmwwWXfbRAATap/kg1eJqJwY6u
DTcidHy3ZD/qxLwnyhHuh2pWhqhTv43ebMfq43C69i7Zts3S1bjoRuErolXq2iaINMVG+GhKU73m
1tmenU4gKMImCpWtELDuVQLGRFcYrzUpou13rTyOgkqmYld+t8S05yHnCcRuECfuxUX9VNz0E8AV
9ruQGXudcqqlPcsX9gequ9G37dYdJhGqhZZlRnFwDSE+HVDTv2JHMQKM356K1o4H08icwtwTicfM
wSAsKTIHVij29EU+8YvwH3Mz1nR4hP9JwDsEHquG7yraAXsn3sAfaBuEwo5UdNVofvI+JoYVAqfj
YqJ4QFAzXJXrGp5aV5MFzB1hMPeDV46FneheukVwxtPyKgjqhfpsfZa8/huZ+CjUY0itPReSubS9
VfFSNa5oJri6FTOqxZuHXzAtJGQoUI/Q1LV/rp9XC0ZYhaEcuWDLm1QlcnJKHv51lmUtTlofMZYa
LLBA9mDv8e8CnoI2JDAfFMAZW2oj+otg+ytcYds/kWHGmZScbiIFQVrQs69rovRm/O368gri2AdI
hyz7rpg7+HPeN1FVzr96tm+OrEy4YvVKZuN7ccwj0sOVUwNCKG7W35qMzpPW+QgRoc9GVb7TatEw
i9V2uHgNeM2J7sYpCkNdX4ppp6uBd6OVqOh0+nTFOFnyZ2mQugkMRrs5PNQ0kdBMNgd+SuKwq9rG
1hz2Lm2ehhSlavx+jfEsg0VE/1G+bjNvv28z7e/wOsNDd+1X3dwQvasddqUVrfQTgSwJOwxE7727
dOHAOdLOh91k4BV1NLmZLDIfezUkUkvEbW0KdVYWhcFzFCFBwEQmpqP4BwfuwjIbJHFEZpLmCgmI
23a9P/nZQh2L3iabA9sL6cmvDuoHEOqJea/mTnrT7zeuW4sOpCDxCMCZG9dSRRGhIDA3dVT1M/7G
G20GMrbaDB8DmtFdNtk84ACp0aqtK5ixnOCY4dKeEvjiv8xfqpgN359JyS8N4bEMlvpNCMVv4+Jj
J3+MryUkVr17ZTKMsB5lxygvTPzoYybhBVztW2GpJKtcZxAzMRfofciq1cO2uT61FNpRnkP7U1YY
aPs1l+bVw2Q8lBQZ7IMa0csQXnBtBCxEeQ3kPFBVVydj8jJSPKSeGNX9Y9Gk9OE3UkSI6wM38qny
bvadNhkSGPwsW1GGNLNF62xh23k4B5MXME3jFEE46f8Y9szq80VeLo3XcnXiFUNEQzkQAfmCJiZg
uXTvMvT5F4mpg9835F9qh7leUaYIT/Drtj1X2pB5t+T0cd0ghnEamWgJNj8KVGzOFpo5DQaWoCMf
I8/K80Mawwip7dQIa5RtxEYSPJDqBt3Wn4YZOCGlIbnv98Y7EFZ6H5C/gz/zEfjU/Fgdf6qD4FU4
K2kvZkcT/4DE05NWJc3HDwWuthSRPCF3xojvki02xT+MSPLxbKw/poQo4jBPz8h0i9N7GeHaTMJH
h5n4SEGPX9t4r/H6HGcShr+TNpzLS+gWhcYVmK5bOxgtAxKN0iHdHz6GyfT3AqfmdghRwD/Z7Dkh
MSbd8huILED50tE/wOFzH6TzwLdgu81u5L0SknCwD9eIkLxjYTEiaiavpzxvWMlvqdKbJ42h8UiO
3ktkVmuPHTJhMvM7/T4qRA+6UiPL7k9tpFIEtC9QojoX8u2kZg1OZEiQFXs0WscaQA1Asebw1ZgA
CBuVFMj07HTkttrDx3iZFWBT9lE2sggq+zbJEXFl+r7o3XVJ5kcOBy+8LjOJHjSXefsv6ye0sZxV
SOLRFj06cSsLAL/m7VtKLUD9WocukipMCH/3EZbZKcN0k0Gsy9LpxUmCbjEaTLwQMof6AsFtqwXB
E3mpcAMPZc4mS8nXbkSYNzJMj73DvtjJnpZFhLDN29NJJuI5GgveWWpqwrAirh1x+LNVQyZMN6KU
td1FfJXgJGdvo1KpKXzvxsI3bNDaLBUXVpqDqXMHIc717gbjKNPUDG3cAxv0SoVPoFBOTrkxGmUL
ZJi0DXY88mfyETLFXNOWZr8GddZNmsFn/5+ctCGV4a0lRQkGITIlRKd2nI/pqS+ArLLbT2zxv3gp
7e040YWzmb/ywsvedX574uXBf7J3gtSmMjpmlBtzk0Nit4AMA0/OyBXJp5Y2xySuek7xb0MEEcvl
wQM7MlzfXAA05G3ZggXTo7o2+abcuuWF4i1Ib6yoMh7N2e0Fe1nWOxAnpq2WCO/M7chauvlnCKQt
6uFX9rFcbRzuelMjdlQ25Ts112cKaBja9AgpYVx0GE7/EpI24WNrJO0RL4DUySUU7gL3TI1qVI/t
TKPOl5ibcXTnkSxf39tIxZYvELPUTNO+RnKXAa4Han0/6L6KiskgVHjEK22dAcTfG+lvU/TEpRSw
5mxzeD296zfrMRlJW5bbj8v7jofo7GwdESs9qUrYuQa7qz3Xd1q2WCGzs5I0tqPqyl8M3iwX+RT1
LKZdAmNd2y7gg0xuQe098RVg3LUr3DO3NkplvmHRH/Dg6pjoXTfwVkzC2SrKrhBYtWiKhlefOEni
H9apNUYpnCnH02TrauIy7EruuhrqM5/qi7RZbHYDm1bvYQ9X6+y8JVK6CnrfS1RJzG65TE0sLHj7
lBsalur+wmVCir4Uj5O8Z4SVg2k44zkwZoyYf4N8FxsWga/9tXSG7rb4Et5Sguujt+jCUhGh4w0u
D+wB+OLirNjU3PD+o8PJ1LrGu7u5q5KWjIXqCJuJ6wA4XG1mZtL1XgHC0a/END8xwBdGoM9O7HMK
kfz7M6K9yPZYDRHW6YrDIk1hx4U5wIpKEy+90UysuZGunog/1/RHtlNZm43OJF3GRnZLXRcNHcB1
iajN2mytoQBvXwohqm0rHnxMAM2tNFjQhBgNzDEg+UNhtwn/xTmI7v/HtjEosrOjY2WCDsbPhZDZ
MDZXTCtxlzI8LZ7mNDXgYzsLRea/UKwBMa8F7Y5LJ8ehX3HC1MCT9vM4xoDXg3LrdUdIE3NiTdRD
hOME1MMCE9CVo1LM5lo7aaHoE3Jw6cRPasFdqTrUa5g+yMGgSTHRkT3fix3O1JENVmahdtRClTNB
UoryI4Iy1IwZHpGLbUDRCg8EiATTndMqaneRZjBXzFsRxaJyNlvNOuNfHPJ3uBHCwG8rgN/xYV69
Fc2fQtR2Uwt2LA3lBUHd4sQ9EbX2kJUwVerRrA5q1La3FcTepa3AK6aFNYz7Y1+S8Iw05wLoK1O6
tKAs+bKTVYctkpPwxnESGqTVYEmCEL4Cv+HA15vAmiKsG/CCWJk8iLLJx4t7tkzBfSoSk0L24lD/
qTB81qn3yCs+5qST1fJatNdvvoWQGhftEysJxzs0ju105adIdH7pUePRuvW2Ba0wypLpZElMJO7L
j24NEmUcCnaRTC/BXXF+Mz6lkY4gcOvQdgIaAUoXiG9ZgDl+oIRaxC3Ziewn8YgTMiEhuEaOFyo2
B3e1apEHN+cD/YoxBsJW/o6wvYkoE7PTsfWZu+2mJhtT6X+EnZqCSstZaVplyULXNIXSYtoL0qIJ
sm1ecRZaKiRCa5cDTmLE16spjy55qvqPFBkL8vaoEeJFEschlnwtXJ+RFRQFjg8SKhEfINyBwj3l
f6erSQXTYM4M3B3fv/ejg0RguAHhfCAxJ2KQ1NLw7etNjILD80TjvnzylSXSyE9d8rz39ou6YT9f
u5/RGop/nZXf7TbzQsmkkoVa04oCML3mMYEGISm+8AGkNgjOvJOLk0vOGILYsXF1lnK6AxnOYYJz
4I6jc5tTx3kUQ4/uhE4qe7TxJbTIjZnulYEDmCSVrsOnSRkngdEDxPxnnLmJY16YqD0b44zih5dx
JPY0rb/oC8L+E1gt7cMnqLsxGkmIA3GCi0TyUjY8fRD1IgG6e88a2/fn18t0C+pAkHG7RUf0Brgb
AhlOduGfFEVvA2gZgZnJsYptW0yIgLZ9BDoAWFlF3xZAKkoFP2gvsHtXTM6KXYda0rH/KXeoKUy1
NF258/YmnuDlfIypVdenDQZfU9/K/22P1tXixGxoJddZTJ+JEHIoqAypAR7NxcJ2riBslwT2AlHl
prnteHZWS5wrGNAq8w3Z9vZW8xawljnYh38ahqU6ZBk2udhF2T0p/odAZRXLWTlD++r63zJMnOzt
S03yCQkWK5B/VUgIpfdijHYT/0yrGUPWdzKuwyBMzZyf/a/Jbqe+AJ6AyYUM0TOipbAv0uuzDleh
mOBISoLxrry+daGrHzEo8bky6iPTx0TzY/wZ4RJkHwA++lfjKYGkd1W1rFn1RcwPqyxFKHJl4SFZ
2IG2Jj2gn9fvQ1FA1G58HqvAgGPAqhbqw7GiCrN4mB3zFWNVoEHHXL3B68u80PMEwfLa8nhc1beP
ByIPgo+p0o80NHZ/mPt2L04Ut/NNRVghQG+YB+R/sqvCX4ZIpqmvpJB84CcEODFk37osIWrROSbH
JUokjRk8M7N8/vVLWUYmmO5bXrtLDG/9cVcHax/uvY3DOITrET09SBWzW4vIPaAD31rsEVgBvbVN
OWeIJNcthWnc7OP6q/PZhH2Fs0sSHrM4Xfhnjdih63UNPdDEDSBYFYMAxuAT3t8M0QsVHcCpkrsv
KeY90CoRCE3a0rA3iOqhKEMveMnbb+SgP5oGzHfNaG0BsPb+EVQ2UAiLP6kARp42Z0ajxcGJtQg8
1QCiI2uPcIL2LvlNo4qs++WUIPYbNyTPpQyRZmlDf0LgP36mMYbow/Dx+ywLypSiv8m/dbJGLK/W
C1i+CGDiTn/8wmKu9puo57Jyw0jG2NZRDZH4slrymFbuqJbzOINZugHlCsZbIlaM/qz6B8XaAibb
gDtBVJnkfZeXrCenusaaPgsRF+m8UIIMOtK/U9mSz/jFGORee3kzkNkGjY5xBSXx0upkdlbCAgGy
mwNy9JwFcG0mHqsoC3Q797HVtd2HNooWbmzXzeW5Dmm2DuT4xdYCcl6j/ltjGBfGLMCi+DKgp4Os
dLjjx7BaphkdSKTojEEfFE/oIRFyOPtb1KQioh/9fUf1hl0qKwUzxNXS/POadKIOqvLwXDLycdhH
RE8rxoWK1zq59oI+M26WveWZTOmHfzyco81naOIVc72FAJO/RiyO8a9lkwnBtYjzlZpRiAKcw5Fo
+Sxuxxxb3y8eMMrAAgV7qpolJNkcH7WRmtrgLwk9gS6uU+5SLywPtTsGUuVU12KmK37DIz8Nde7U
jkKZ8lbUd5GrcUHdYOKq/LEu6Y9Cf6bzkfthEUJSgFlW4A05DA5GrJKuJ78AfPM/WkjSMc2HZtRC
3SuddHe+rtqOiAbvZx3NKeypAYkec6qfeAiHOsjJQQlW/9UTbYg71Yns/50B8zaEuLlcjAAhzAZ+
ykV5dmZd2s/hAzegsTKtXUcXm3j67WB2qUFejlG0ZYdNDe4Q+xa3/GF2LuWuj8ClDaLY78/hDJrJ
PjRQsKMWQpmRsCHh60mvofbPl9PsXM3BOUq6qUg7+IPEC+WE4+xxwIQwzVv90Nv1xQxnDIJZqsXK
VFfw9zgYiDRrmyKhtY9aJL0yjFE9TMvBl9C1OnNylWZBaaIGj+G6OTMOmdJe+ujO0TAg99tDVUIS
lC5cbggLzlYyHyhS8bdsyAK+2bX9YYzmL46Nc+DIf9zbYfg0xYyliVn2cGxNf8Ro/az7cvjLtRvm
r9TE9kxKnhKmlnq3PO1t61HU05JSGS4knMlaTDOX8mJ4hlix2U3v3pc4PijhFYA475KEidls/SpG
IEPSB5OTN5No6GRmsxW3koh9E3HIzpdAJPtw3BHowHJ44ADNDrJn1FXj7duQdb703pr2vdhIfyV2
SaWM2POhn3n8hTle4SPCZXy03pw+9F4E0avOWLkDI8BIRo2Nu/58F/Ax+bDmV4vmjgAi92jCQIge
JxRuTd+zX44QfZl8CB+toX7Z4orjqw20ft4LjQQLp4gdyxjnOWCc2R0wVlaJpQcbFSQDiEmsxPkA
JZljDkDIXYT+NgfmIa+vBOg/7B2QFv1gamufFWQ6Iq9kNjTTEpCjr5kADhFepwDkdxmEe75lYLj1
d+KqsQJypTYoGMwrL0wDi8zlYzR3ZUv9WPhJnBNc8bWX3RhQrzWJYJFt0rRnfcOsTTznDmqK9ac3
hTQ2CO+bxoOLe+fOMG9w3q0HmjI9dYPqPHqSnfIyfAZio/zlrvErdIrXgxTRbyxHmLKXFHoGgQ2g
kiL4kUmOpTfnhqzGsduxRLtP/8Vrq0T/WEpZJqXFdYPiFhlvuvDGZL8J6luA2lK7M8Yy1eJ1hWzY
2KJ5GHZqdo2KVl65jKVzESI/jipZOUAwANc+FlGWntIAKRsFBNCXM2uG8Ozg+/uGPtVreCIxKMkN
+vjlgz2Wy485y22x0XkPNwqLwb2dx9qI+enJ/oF3NoelSo+ksIcP8FCyZ255pcWlU9QZFt5Pu5R7
ZzoyLHWES+RadTYsZk2ePAdybyzOwgj5dMAH5Wg2bWrTJIg7TwoSLlya254XVs7wiIUgYbd7vFmG
8U0Pu2CdoStR4foq90OXXrGkkCeYuVCXPTHzODFX5MLeXDKoV/pag0J5624RwL4NgW5MGYvrk6M1
00BzQYaeUCG7IUBBG/+aNmBMU5u1DsPlPbRnnYJz9HyV0/Vd7xNBxx+G6eMJV6/7Q1ctV2QYi56a
hC18CTgj4BkcpEI9jQILD9g/csN8aBM6nSLz/x6RDTdrPINobd8kT5OoS4UHjmlq5qe2dKEuW1ah
4duB+OZi0rF886mC6ELm9wQu1phPiJckVwLjoK2MrcFUCvsai5FzaGicUiKB182vvbDhu6xgOcnf
UKwoKD33qjrT/Pyyc9rmX7UttjtTnjSNPZqrrLdjUb2CO1cIdJBCK7pReuotMlkbz/050HafYddu
69APIKzc2IF2KkfNOhRrvirHrJHR8F/kLYy3ScHc1DZnnDU9UIxi28FN8t/nxkhjh+h+p6gh4RVx
939Vt+nG40N4Gyh+LQ6Yg1VWVBM2+4jHAHYM1aXm5fQG/nLKVXeKTGZRSnv8ifReD5HSvnWynJUi
6FOQ5nVp0J0uYxS9T88+duV7qasGsQKE6noGqFuxKzaYO8HuHjYMuKD59tBo50/4JWRYMPanFYAG
efEgQNRNw+2d134IUIqbKxU0St4wDGlE5420pPNuQtgq/9d94KggWvKBEw9BVdFNlzLGgIxTGkcG
BdVln2yYrD5IKz7Cf8/j00CKCI88FA9rOeaMEzTyT82ORewQU2v5l/ltZyXFNY+nSjc1Rw9yixWC
/N9Y9z4z+O8VXBuBjAN61bz1l+0xiItrajxureIhR0/AI3xOXhTnVRmmAx38VwXkx1qZFDog/oG0
x5COVVGNhtYORVHchqsEisC3dkK1Q383bOM15lYvInp4XJsXN8IXOILac2XBy9ko+aBR2J0oMWoB
XRdwDWO90Yerkq1pBUHaFc4YHIqgf6BevXmCZu1ESltdWNb2J5iqHU6g0UJ2rCpvNo43nKYA5SyR
GuROIBXXf8R8rtq8vHCGTIZfkZ49n/LLnTg31dAfZ1kUCJyUjnAK3k4JKtSU+G21pAp/eC+cuRvx
qdAy6ImtflL2QAUdgWAO11vmjsT6CAs0fs68lIIaYGY4JHQfANO0BZltkfueLiQA9UJcbyOTJaF+
v0AOnHkf3DO5EYPp1vodzdYAve6pIPczDNkyzjUpispyunRSOxyAqxxatYwcD+QcS9zV4qH+biHO
RYqJsTFR+LAzS4jmWUY1OL33zJMyIIp4KLwDMcc3NKtxAPK5+rTh6grZTmhRwUazTHIQHLocHSz0
BtBQMyUuIlOMHjN7Aepaq1YnY1diRxsUctnPp3eu4cPMnh6aROk3pDWbQX/1ylPEF7pgFOPj9Fv/
ZbqeTbIaYrovFFuXEkHvLnUNaA5UFKMIyEdoocme6BaLdUCrgkZ8zd1LvYQBVQm4LrcLlkErrLDn
cT8zBYnu8JAWOLRTwEFkFPXs5qn9ck0qwcX8oBg5qF83BS+mvHAulhC5Y9EgnPyeH46G97jOCfha
0mHMXB7QNPd2sbntQT+GS9TI43smM8RcdqOCNwajwFLFmP5q9A4BjlNa/RnwdYYQfTB2dTDsbhEX
Iiuk4pcbDiQA6QmKT4cpLCYUufn4nxkvdEgGWmIHhblbaI3elNF9Mu+69p1ClyGmsXD1VSbG+SII
Ixx7oZRE3FzeYJgXyWQ4F0Oi0SysGUFClDDGnJQf1iRZkDBfCiDm68bpaw+nO94PM4C0/I9hyCtC
OKrE4yWHlP85nAZ52OSUX2XKCy5dqgA5CdnOwK3lZl1fm2+JyMoNxnVt9vD6HQGVwlS6HjH0RUBu
v0ZGClr/rlvf47vQW/sRCVeo/IW1+hgKZxPMTwp7dFKQhwuDtSgWOQ3hkugWQHZs18RbFEn/T7CN
jaV1CKeMtwVeq88/VBCM1b3XUu8WhNMnqDVI37ibpZvrKL8cHmrMzfiTEDHzvXp4PfDDceOlFzE3
DXd0UkW+L3hfUvbloDBXKJPURZsVdwyHMXNYwcv6zM0xDyAEAqw5Vqy8k9dcUQSEjDZiadW0WXJW
5VIhh4qqCEzdy6+BQODKkyxMOkGB244axu7u+HQyAgs9UNhytu0nqA6slSzTChw8UjRWwXDjABwJ
n62WSFpKVBZkZ61j/kf+HBrQ0lY0Zu9CLyBAtUphobAAPgTGMFKrr+SC77jwUqzoonSoA9CLl2Zt
ErlJ2YnFl6Tq4SUhiBy7keeuLH/rE6HpavecLZ61FBkuJDgRjgDolqPuZjmX6wymFAoOM9fxFQf9
m0Han8ebHSafX3rV+7apNU5ForwJpDz5IQirjss6jSaxFGnqErk5EEZf7E86XXLGCm4ttHBi3dhD
FuKD4ADxjMnAa0zG1F5h0QygflRMfBVJMW4LxoyFZVx1nE2Ae8ZWPrN8sC3iw9mjYwzEF6tqB8cL
dTAFHNzhPzZ20HMX0mK0qcqfbu3whbsQQX4W0rBirm3r+PJ5M6IiQMJX/Ep4Te3TTs6RH2lha/sT
01MsiV+IIlqol0HGhginpsYVi7RCu6PNpDtTzFf3PHjqLTQb5W64OAcLAK0PEsF9l5jjZsh1ZYk+
Pzxycxvqnbn25X/rxrrVZNtMTpNPQtSo+sISxYZb1eFCv3Jp3FyHdDKpqmG/IxJBmBTTAA1xjZWO
bXMF/+Zbfh8FONYP10LEcwiLvjqM/TW1lNu7LZZ5MXBJG3SCcxj9ruu8nqGwqm1aK4R4HYvOs0Sg
Wb9pAxO2jZpbOV7k/DS+uz14m7IqMJHG/gvpkNwKxdAG0IdC0nGYOVzahB6OIuSVbTkqIFzsN/AR
VWOf9IC6yV8xius/3S9QdiP0UXav2ENwhYI2DQGEFzHS/KR5PQyWTsDKdYKbdToFoslYx1aYkP4N
hQiR31+EDVfzubfxEpKX8RvwWMPb1AuFMabwi69pRXCG9o+c+8L8YKIM9IthSLOl+LdEaT5Bjl9v
ywPE0yN6Y3zn3QMMxMu6RAF4rBKxMFmWeIswF0/A7k9JwM1exlhAyjdCuRRv7A8CQ9mg6R/zfW7y
vo8LcdxQIBCvZwbmQ/6NGjpbcJIHvlwB566g/74KLAL0h7rAqiwtLkTYZDs8MLei2BwFP8pzHPSJ
8ZgdXScBbZsVC2JgxKvYo/FGkcd7ujmZwuVW6CaOWCMIbGRDOED269VJI+PdWY9NyQhuCPy6G4hz
iU2L5YT5bg6NWwcXwPownuJHHiGyzLwUu2+WqBGcEXz7vK+QuoO9/08FUyDk952D8pJIQ2LFm1za
hDmX9r+pU2mb/ekAUPnaccT1P/TVUaHP2iDzMHA28lngqt3Dk3hHMg5Y64AygL98I9thRdS+e4R8
jBpFVcBwBDbn5edApPZh/w3TqIvB9goBBIZmUlHJcoSaO+XoBxI4lAZecMbGSssy0I94neS6ym2P
tm3gH27DndRuyWNgtqQ/i0lhxp4hBM1JzIztEcDT/vUkmOUIJDUxbl7KKYfHoFW2AgZVRVcxOnR6
fC4xIl6/aFAnpSHqj0Mt1TpN1xYKmLjI2t6heylrRCDuFEb0ugoFw0ZWCRqqaMAD91VkKwMG+i0X
6rkIPdceyEU4Q35ezD/imFKFZNWaHByt4nS+/9GO8lelK7UeSGu3EA6r5DKR+YK45a4adR3YpUAq
piM9vS3PW/TyXDbyoCRNaDIVRlRDCkHUtWo3UaQk7GxcTo+BisNcHnXX5b8zFJhXItxVlcq/f1c2
PYSmiz1i7ixq8dKzLJWt8m8W+dyUGuy/nulhC1uD/CPJs7UrS3Mta31CyJ7blflvcqbWncq1U+6q
e1vIN5Rgv+ormdAwsMrN4Ny9s3SDb9gihY7qKsqUjlR1xVL9G1rDWNAcDPS21enQ7zfg4UBxo0I+
83bQg9H+T7SYhK23dlFosFMXvRjlqOB+NWyznR4dPCN4ijUKOGFq4Gk4xxVdmWtm6yAgk1U9RC+m
n8/hsf25a4/NfiXuyeMdpY1r768vP8RleapZzRxm4tBoApseBomFjFtRvdsG4drzwQHif+cNl/S1
GymlMZKizIrglSlMoCcAPAI9JpPihv0zpTL8n4YtPeHIfQiWCUovROUjOjfukUR9+lYVt7KVavg8
OleCk1q4Ef0sAZh6CddFdkKZ18ZtqfRJfXH3os5e5+g8XmCaj5DgzDZP2gCJlbIg26WttSb+VT4B
HJAFoSOij4i/HrBKFBEy1O8INRbBbuoFashfceFEzF0YTrYXU5q/Z1yZ5js81sSYBnT4vsulfNGO
/x79fXYYZmQdgU3l6rQjrPdleX1Jab5SJDGtNObhCQhUMoYowy1vtEZxgUAxV/Gw7fbCINhakYOO
bxS7y8hyqsxvn9pm4ZJVqryn5G5CeEYVf7G+oueCyF97bYkJ/zGaugMRUwks3zs2fTh+d10c7dom
KxzKmhSLTx7pcaW7YwXv5Y6dbhuFdGmftCz7A8H1TbdMKfuj407pJDB7JpjHLjvgFW5vOdCRVBuC
Zp+a+naGB44D2pa/8Y2uZpaVfDecfWhdPwpfbeiFSJzhgO61h6ku9Mb102TVp/X3U7nrtaJCZps5
LXiFwbeFGdopBvpsCpX1IWOkQn5JeSHq8wVuc+Rqh5S+MtV64Bkd2rDWI8OgNcdQ1QNGKjN5Gt9e
4yRlb7GbyaGgbVGGEz5dAlADpzoU2PsEMT2shFA88mGyH96eX/ev7NM9YiXZIMJ2a7AcNsv8tpp8
qfGThU/8cNJ858xnxST0ZNS5QHLEt/R/G3dNTmHO64AOBoLLUAHfTpFg5wkRTGVrRHStijwl/TbY
vJ05EzW11/od/Ug0gngRnOGruOx3e6CtsYgtZ/miFEK7F0QeLUnr/fOfLLn3CflMzOQeoaGMQSB0
/OcTS+boAwsAzG7EX6JgwR1IqwykN+xE1fpdFfoPNK6X5FJXbXjh9uwHaEYGynuFdXMILx/J0YGN
MVbE6HagejS7bydzuKu+fhNrcEvuHUvCLhpKyV9KucY7UVL+P7hvSMW8OjU7kz1bCzkNrDcqC5g1
H9kQVn2XmECSvRNFwQpImOVk8kN/Jb1JuSlnymmWmJz7tNiCOf0CA+CE0pMBtsn2qBfcJwPYyEYk
RnAoXxVWBEKCTCvBoaQDzmKDHuTy0cgZyzbu00mu6HgD8GKztqy3vx3BU4alqRLiEpRBD42+Djz4
/UEUTRU7U6hYFu2jvStmxGp6rV2PHPJalpBUpuJzd47URUojve3WA7J2Dy884PWv7MOtJNmB7ZzI
CfYhwRBUk+lAICM9vunnKSmDwECLT6OAof87Oa2LJdJxw6P+d2lYXqytBY1EzrfXRyw5f2UWCSN4
xp3BEApKN9/8Jd6u4bwT42FtzKgCWm1UudaxOvVDn5Dv5HmnOqpCXMNb0QhAtygX4YTrYJTFACIw
5EjZrmtzjbx1XHrz88K+NykwTcjs+aqRnTGwXXihRnCEMPyKG3mUY3hK1BEYFN4/edqi33UXkffq
2HEbTHUjzB7UxRfKUHngWUM0f5j45eZUcSGya8UlZG2jbRkdai3Usv7e3yd27ua4q5gyNQ1qo2+m
WCj/g0jSPy/hxb0IjGTZx+tjvzZk6UxHEOJjNrlsCWAE5a1PM+nkGhib+KlrR9cs6bIi0bz+2y4c
TyuJD9YG8Yu3Q6U3GIFoZGGOkK+tZN90wTRoQkLFz7j4Q5pmHSscbW+QGWzGXfeaV+5cGUDvcVXm
CP8VTkD1HrcRzYhK7uOg2oc97YqEi4dpuTj4eVu8zzKQMVWAIkwZKaPgWuryVu77djxmZ6VVCqaa
PJhvWIehU/8PlIrqMNiL1HnVaM+yqVhAd+CYs+t4eHUmjSgC6EhSRAp9cHDanVL/yeORr6QgObs8
J5d043RjyKeDGBnnQxzGWRbaZmsKoO/Hu6iEXsmfR6zin09QA58RwfjNeAVqlbwvNuANMHeZmJNO
WWgtSziMqU+Kqur/lKBZypFrctcG24l9r48K5txLvBWRcSfr3qkKu9+fhI3QqAlgaLYRpc6XWmEN
AFT2oMZ/cem5VLZ/hp753o7xjoOVNDZsNSoDB+ziKIGyCWIglEoaGpGQdvcxTz5hApxUFksZTVt5
4RVLz2ebJqgSE1PApti8QWEcXgOfmUiGU8uclyN6Q0kj6I/dBLk95phyx1Q7uBBVP49w9IVKzmdM
jour8MEBVkSvn/9mC2hbDGjSpjCtdT7TxwwSTgq+vYp7A3SsQboRqM7Te7HlQLY3x6KnwqwAdm6Q
mo0ZUqi//EqzZtek3hxKH9LXmPgQ0iqNS6QLnRWqLRiynXs/wSr3XqqpkyicWz2CFS4tclq8g5ds
4F6yd4qrRCegllYQQDnEwgMiLwP3A1Xcr+bYlPuxMgFZaZ5STkoqPV46eu3aSYRaP/x6cVHDb93y
4W8GT17CUQoWoFLwoe+FM93bz1VPA+jLZchfIvzcOXSGvNL51G9FcgNONaaRGozSiFzJJQGJtead
pqDvC3wjTbm6R9gCSpX/uP12IBIMikBcCOk+yIejLUgwYE2GTaDPQXy6dVV3mXCeX4LVtf3dgKJF
qpmkGZdk2OyQcYEggRHzReBj/LDOb9i7ct+FJUGq7Rf5xKtnfG9RThnrLm9mO0yhUpRfTcAUEwz/
nJkZHW+RJrmWcY2gco+/mskA1iNHJKUx+5UTa6WUKroxs4qidADbsrGzBnkeK0+lAACG3brnfs/I
1HE3GAprY7H8anvuTOuRshD4Hiv7AeHytWzU0GKm9jsx+2GWCYTs4I2P80bv5Lt8VbA2hQPtTUQ1
ur7hAy6B3EIGC6Q4/WXUjJGUMjHPkwQx6fWbF8sHgD4G9BJd4lVLDEOzv6jTRAGs0yRYJlwvj9x4
JjxKqv6Q6FMxdOd58IbORmqknR0ccn4Nv9Og5k6SHc6Jb5q0MJJRc3l2Iky00PwrB3sHp6gfvwHm
RkBWDBfxHu7aaaXNLXJRvkB4J7pRH0OZI0MC7w2ESDHdChpfAJcur5ohT2LD+FmfBl7HrVFWkuj8
t2z7i7matfRTCiundQ4EAmPA+4lLaTV1qdCgmbK5jxfAoGdwkUz7pGR5TD3bLSqNZ/76lQZMMEQM
AzB272j/JWzmUQa+Ls2wEwBPao1tBycIXP+hysFKzghwP54ewu3zJl2tqRBDrbbI0xjOz3+ec8L9
tWyLgGitDSBKA/U92b4UvtQURI3CwQ995+X7+1F7ZYhI0s6K73uJSfE6QTxEoTFguDHLfRoFmin6
GI0I2sKBSfcqdw67zimehxt4l5rFMI9Wc3cue+t5Uc3EvOgttXAhauREOlBSbp7uj7LjSI9gIeIN
+xg7JfkSFqJIlDehjOjCfvpoS4BmWBFH5ckNUTC1Pk1LuyRue2MGth6FsXtBZogDNAZ6s4mA7yYA
LJstALIb4DvTSLA+vFshVib76CyWEBGeQEgvygbEZ8tcFD0Qq8JHBK7oxYQWWzZznmridytVetvU
dIukBY4wyfK/jwBWzYK8MxGxOrmQWSKDM+X9esb65NC6xQTQsUrRq5rl6KXlakPBZRiW24utX8fp
wNlVzXNkSz2icdlIzJG+QTrM4hGvh2HiV1GFZFmeFrbM/+RFZlJEb/rpxN0R+AIZavjL6yKgwNFR
YbUCleaaWSYqV6gzblt5CFV0QirmY4GIdLJtCmuThaxkX6U1P8c/QA//nx1XNzMQ3JCGQQ+l4i/z
iVYqg3Cjnb31K/1yKhU7Ck8tcP1DNXJjdQSmk6zcgTsS0aZSAiwLkamcuEK6ufyhZ/GaO+U8vWYo
q/GXyxl1ydYtvEU3DzM8L0Sk0dzP04Q8KN0API0nz1ZJEqEuBKcpbDEPGcY65SwcoG+HhpekHRv9
qsq5urFK/jcovrhQgeFMXGNR8W8M4d8/lXcw2LnzY0PrjWpo5fuGkioiQXK1glNGh//47QJ0kEe5
dSVEgpHz1qSnbwGkZENB5fivpseYh8nyxOj+z4TT3/QqQJJgBHA8E0ADle9oWqKY/3pHimHvi5v4
ovSjNk4nkBeU7eaxEk7It/TTnB/w+VCdYNidDL05qEkFoQTjU9RHfJQmGjZ4azluCgqMHTCaqI2+
0q+NYTC8nZdyOn4ZfcM+v4fY0TxMIpn5WRvngjSKtUcul4g6DGh8PVly/APs9I9myilIXIHMn1cF
zfzDGRNPgtP6iHQSo47G3mQUnx5PeFSXQsY8wVzmhxEvSPSR+lAMZ9G0lyF8lToNZ9re8tLHZ2YY
CkQ+bH0QoF++Xvp9rA8wW3GR2TA+Y2rlany0rrNJdLt5KTq2FaDrzXaE4KwJGU4/5p6Prl7W7e2A
TMrJjgZtFWXRqAxywsHld9ToT0C+pJBzyNrH6ZyTmNIxxFi9BeG5W/qHK1G56QF8ECMySA2INqQC
uKViEskIQykmVOeyHlnF2ccioSBSNH0v6zKEvV2EdDz+dgQ8WxuXVKwR9bIw7JFkKkE8BELSYL/Q
mss0SSDjBZQICVO8bSn2QJSeKhfaeo9pRpzC1SnzFDrAHNlkQWX1XevXIXGZYy06d3UeY8Peb6Ns
FpWDNc63BCwIZWFVFGfgdkBSAH+wH9w+XcqyI3zK/41BIJcwTKg9uNJZOPjBCAIvgwdUI3tAiym2
wc1LunO4SfqfFEcb9LYZreRELCDZiIt2KU0VzyXWfy/GdLuFqw0D9AlNYKSAVzbrvJ53oJXiEPDz
Y47lGbn4wFu7J6xt7iaqasWYeWFIOXyvISsyj3NCNa3mOB4HtJhDPMV6vSdWApoLayiJXuKIn95N
OPt/ct5sBiFyiKbx4/rqqftXaLcVvyKYRyI4mPmWpkooKaFCMzCNbSZF3RicsdAKeQob0IGmJEHJ
HzFSplG8Iql4RRao3SLolTUAVwPk/62oSS44dnnt4gNrmw6Cbv0bO+5GxDDEDEp9gvhUm5skfYy/
P54XSze5lr+TbQ1GfhjWDxeu7abEanf2kxwNw7xgP0awVrxosFdvsVvUVPsueesRyAGOHBIQdLMo
kXo2BX85GL4VdWkN8NT0CE8t8tLmWMqi7VSDquUFrglaqlBW6pjipIqcZPNpO6kV3CZbauO6dYud
w82lMze+sUN6WILtapE870THAMR52/s8VPYqCJYBjiejLWBhiN88TE9YL5yPwf/s363tcruM+4wi
YClY0CaztZyxH0E9s8P6BSQhIPrCK7ROSRh6+fYgRvEPpO0zywUgKB3MGlZ73k91CNDubLDMlVuM
vLh5lFHWrLt5P2DiJl8m5ZoN+XEcymDsU4k6wViVOV3ZmnSBwCXML9NvqHdNXlFgKXBk/4cLWgUL
A5tDH8TGJHQYub8xtlJ3YYj80w1fy/OUlIuSJ80ffvO/rNJSjHxAvrbF9r5YfJH5iU5of/Q4qba6
v0YtvRzRDx4sNdG1dBj3HctKyC9R+qe0HuMY6vmbDs4k9FfmzJ2eCOkLAeV9aID0bmzg/pP4r4tj
AkBtqVoQ73pFkre4wXdTckA1/1qqSKm06ly6tm2QtGXb7vmh+xnbDqnoQS1pBfLMlX+IyPxZ3S/B
TH3i0/d+0rgJfn8abodstvgfTLuFOgSJALzZZiwDd60EhZFaTr1B03DfKGUzpeAsa8hW74A2WlvM
NUG3qfmPj/9cLnnNIt7bTc8rPYAz1vGsdMcHmwEXiOhpX7YDLMWuDays2x1ovxyeD+6ITXXU6Iom
Q79LCvbs6knYKKQHO0eRAK6FC6O8RRgvAU6PTInC3P8Pdfj+uMcC3GW4LsJ0rwLlrM/Vtcz1AW9L
fnXQO3RPIIgUWRF57SdtP1EffsbsxNvL7+I7U8HAPIUAF2WRz+UvdFX4JeHW0o9E4Jqw931c/yAf
eBLB4lpddnLn4hn0aufsEnlNpLC/wIckkYW2yfXnorCsAp7B6sSKAJaca5OUUujluaH+ubTDuSVP
dLHRtnXK6EYYaLrtZbscoyscoHUFgIIavo3o4AtiEWtVacJdLj4ix/1DKpVqS4iNe2LEe/kl8bgl
a06CAyCPYJH1yxape/Vavo7IeSpp94t6ezF55Qw1tTjIb7yWgWmd8ktdZdzVM3H/W/Od0FABdPnQ
GjXxt6Y/ZyqNx2Q9/9QrrO7yGbZUpFZkKna1wn4JgNtHiAWMAyaaC/I5WOSPAMrnC7Gcl94JRGog
U00zqkix6y69/ukKjfPsz/P9WbXa7IBOxF6rknS9Ah20rgIpYHwcokU7V+/pr/AVc7HU0xOE+60j
PnrZoGg/JjADFQb7jVM9wTqFTA74JZdI0NNLcejQNt7Il2ROSh6qI52JvS9XWLbHw0ObYYAucs5Y
XAsdCdneEC08OESiAOyvgDKINCSR4EUzKTL1rldJEsfxo15A+sW+Sg4FIZpfTJdCKmIPUnoTag+j
onof9/zEN06twoZKD38jH1l4Re8oXeLadcANqB5xh9bieu67ddjlPF0XscABmIogcbiQGiNSvyfK
J/Iu4RbuqXGQSGBpXfYzK46lV1Cxvtc+6MgqmuvEchpvMsfj4L0YKEi0p/afdmSlpyc8bssJ/C3O
GwYq0fBHiZkkC8rbzvn8lAl3bjKSYDjmHijvDRrUtqYC9/P6/piDHXR32oa3iJyWmtkp4hyg65s7
SDReqBDmnB4l1DZrFdtT57GI3p7ZMhUV+Ny9GhNNzhGlYWSEMc9goqx11buiTXXPk0euqLVm71Bf
K98fuGKJxXBhL4eMqSqucPEmKf421aD9O79vTJIbeJ6oJym6ECc4DRN1O/k64dZBKjodiYI8OqbX
X0W0CSDfWNxpiBk46joUnJsz2AXnEOkOmuf3VypzEHdxNiu/+dIK5alWOr/LB1q101xZB8RNApgF
qHYuz2JneKZrsMN0jjpqzi4AAs4cEcTDoR6hICt2jzXEZkJ/m9JnTC9/BpAQp9biPqw/TPWftxE0
ScbGn56PuAEILfpsTLv36YJWGdZOnWRmKHvR2eP6tSk1EvLxTEa54WkQJFqpsrc9AHxwceqMPGrz
4jmoFNpXCKv/fgosPhViyn3OjA629Aac0ebnW3EenEMIdZFjacOKxF/a5KFKCqy34RkzmE/ZuanY
vlBRtq2cSkRKeYwbWT34GtUyAswFleZ4BefX3PpnU8NEaOzghiN2f8xoXt64ICtkYu16V8M838HC
NCSq2aBj6SjpTwVjK85b5ASf297g3lsfUaBhuEPqAKjvPvSTKNYJ8AIOuUsnxN+Mc4obEfS7z8Wv
5a3symheECD6j1+2VAbe30SPgDOVVXZhZH5H17LiihrvZI2La9qN2Na6LqYBgCX2TmZnYcJ2XbJU
leEtARyEmO9k9pIz4AwFYPEybu59dOw/+PmTBXhXcJ0V31pbpjf7WCg0M7aBTGouqEVwQbMdHdN7
er00RRFeFiYNaNqqGcYpRjLBlAkdKEnO9gMM9fo8tzsuAivM+2qIIoU76yRQ+47pVrZ0fTsrQKBd
EdHVayv4rWZgm8rfFUbT3wuGJJw5aG5uG9mkxR//qGVjxm0g+0XuRIUPwFG/JWQlu7goju8RI8d6
Cg0i/Tr/hLcBHUjDsfgXJO1S2sNPvmdJlY3uJwM2ZhX/XaA9619eLcK1PqWGz+bNQWbyzq59NXzh
JZUM3C+GEkYtxlTMm1fg6pEU1j46wN4vrweSYwfIMjQDxr0I1bPJm6b//hEApmS/x43Y73myftEp
GnaGscsINgud+13llAOPtvj0Iel1NfZTCE+/+2bxE9jvl2mY3fCeBbHUm6jHiH0BROvXqEJiASb1
x7uXiLVLxvwcxXEve2VDUo3n7n2lDYxsle7NTPnQdfjsJs1BIW1t1HLW7uqlhRBymbvSMoNGP5T2
xiCAfEoQTrkSLILLvgWt4zLJJelVyW3s+GhMaTHv3PkmDI5SyiXftOc453tptSDDdX69cDZ0d1Jq
o3w36gtBjN0X0qrbzHS0pqT/XqtfbNePbv2naJ/hI9qXtZOoEk0a3zHLSequ72QE3/0jg4Xclja5
ZszE5/5eEJQ4vb5ZpN6r2vYiRthC3qAgyCdjkj2PBqscSvdVkMQJEeV5DjQKsMqfCDk5lBhD18DY
LKjbAO41lXGPTt8jXVjKgj+kxrzTyT3rGqiDoVCo3dI0bUG8rBOq0mzE+8/UjoKC+4iANqzigDJ9
AIbc58co/A1+L1dvk8iRQ+nQKHMi87gxNUN//TBtre0elPV0K6kj2kxAN8WoO+Z/MIHr4X3LOKW1
/lF3KjpkMZO9Hn2lLOwcz/T0D7s5E7CCN/hlwtF977HJySqlRZc8Qn0Ox9p+ScZD+JdgCIzPO05f
DKytiThfmOydGU0OTjhZFbIBLFWWpzwgMa6BqQtqk6dpoaXFXcGzwxctGYTI4Qk8uFUe0Mzz4BQD
b9evtOPW0FSbfTOnfkNtoaLXNC02Nmco0AuGwIg6hgi/SVk2K4Ecxvvm2YrpauRGOlEGZCu4J+oq
oIM/cTOwnZJVGDYTFgBXweGWnQQMb6ci1USEftEubpZ6og2Ji9/glW+Kj/FpNLZw5TwqXaSYrrQV
dKIodueWOQxG3pCe1/XejkWWC1LGSld7WiPBzOMpLdlTBrYDqPRGxWQzf4S9W6r9V1S5g6tykkSf
5WRJ5aFvwU6rDkDyWeQdwymFx+lhkiPb33oqMxbrkiIerFmN1AmwNsOZLBzRYXJcyuRZzAKzC8d/
fdLFmzS+4AxQB0hVufrZMU9NcRcZTToKhfEWGRx4pSbPtyI42r73DeS6tKDwPs6FBNgQCK9hFhFt
AtldmegB4/MySXZ1ursosOknhdoFasrDLDm5T4hX1PLORWlzGiTL6o6Qkas+N3MA0gUA7PuRRA3b
KxgBsE1KR9jN7f06ISyQ47UnVjxlks2a4wcfD4BMeHuQwNZpdkmLWMQOcb2MKZcL3hkeGjeJQ+GB
uOE/DT+KLAtK1+OvHjkAPCKhtjhFPXqzCeVT+cijJvliDTK5sbo1oF8BY6ZvZvjsj0PeSt0WGz6F
C4WkuEdf0TPY1pZdrQRhoJBBYJ7uQo5k6rB6eIHE68DCSr9sQguMIONymebphTV5uIHbM3PhT4kv
nEbKCGxiVgPNYaLx6PMbb8E+cavu81kMGkLYP9Y9vYvxTAtkbAhDi4XMd84ElPkgITuR6oAPEyKA
/5uds9NShpLeQiJQwuKBuBPuQuX6Li1zPGGpvSJQv+VgoryNo8RKrXJbynv+EtTwlj7uw9gS8u9i
U1nCDH2qaHMl5ZLxGSNwPhDJ6FD5VAq1TvT7vN9JC8pwgMqPXiVaDFskzUAHPwvmyM/lVQuGH3lk
MWqOCfrQASCBQD9tqIN8i3TghyOwKtRTtIxM+5oO/CHmGIrWmDN0vtzR8GcwvQ+DlEwh865jJCl4
yQQaACjX3pvyMI+XxehUbsammEFzm66NWgoI2DdASB3b/CPuPLlNcRp6sI17k9D7wZ/2wiPnZ2Na
sMyxgA9A8A1yHWsGgKRB3rbOrAkDdhVJyWLZwZUk83J1Zm/JYiLNjBs9rpPnACOM5QqXzL7lssh9
eZjeL4AKLWXrwXEWHfRmPyCH3ldT0W478janTGMyOLja1v8K4aTfOyr4LHgLwQsiZCkfolcIB6+W
jTyadsOD0Gvm2wE3fYtWNpMfnf8nGYTd2mXdjrDLSWeZkZ7IE8vw0AMKonXPoHUM2crYlYxJd0Qt
uoDSHhR2zCCeFdJfkOiuR6kjKZguErh/OxZTD9nvY21bjSCDYgr4CdQdllcxkACJWdA+3qKlbAY/
42eWduI8sndLy8xY5IOQWrv/CF/Ewlt9tkyynsncSgaSH4KUjihg+FWoPr+T7GyQtqrmS6KBNg5I
BY/vCKwKPErtoiethvhYWfDxFwJdYGbFsDf0dIErSPaXnYc9UG/QJoXfs+PNaGl+pFn4xflFoH7V
OHHDfKfKmfYdFEtqiTS84GYGwzbJhyfV6oC1poZQL0AtkEwXno1qsj196JrXNuvYgncwGhHH66KH
OjpndAtfzg1SMOtoU1k0LQfFt8EafN6x0NB2Ok9LWN//wb8/X3vPZyFJMsvfQdoHSsidaiiRkx1s
0OTy61/oKL6NmCPyP59pHtTPLieDPZ76KlA3hGSLsni8ZzoTc0bYxUvHGHBp7sPOROfQwxQ5mMm2
aEifZkd+ECLksPkbVZYEkmVIeixf3F/dUY9lEdKW0YiWbDfrOXsFBMqAOm4VnpzYAH65pqxiVgzy
hL8CuZ10F8GBoVXyAKrwIDr43QqBhaXB8POUpHWdB3/R4wdIAFLoUYhouH/syNJb6sXb0k3RhoR2
2M7Rs2pcY3XLs+ZlCbS0dzkJ/OmIRr5osxgfpSx4wKvHZf7Ozl883ETLc5Ellg+oxrRLrVqTZod/
CURaniq0o/I6DWmRf/rr98txusJRCc8IQxf7fc57jwP6vcfmk1qZBziAIZC/JOMaQl+RHJuzxQA+
R1+0yGbs9yBDhLwfEkESoDveAnXnx4Yt0z4m+OZHtglco1ZXIRcR0JCpx8TN7i9GKOCiffkQbi4P
PDhPrW5v9m+KsPXQoYvR2/5MSIEK01sk9VCS/OnoRq3c9/F9JBtLWcn2lOoCzGLCF/YnrVk9wigQ
el4nrsGNkWEjbOhVv2PKSs75jir0KSOTTCpfTiedIAqsquPxktnwrmuoyRCy34B6swQ4nRYFRLz5
7zPHcratjnv8AvMdog1p0dVZaaqEwapn2Z6zt6S//4zxDkFlYXkoCyvz2/Ur+3ui7TCD9eC0e8vR
+ugvVHPZwW2BeKxfFN2wbzUWa+GnxWHohRjhmWQOHm7zaLfarW/irU6kJ+qqxwb/V/kVmpv9G/FM
iX2zArYvy2Efv+jrVCxm+75+TqZ+0idRpzEMY04SkTh8hEnc1NSe5oxwFplDfYQnAZHEH/bQBeLf
mLo2lcwsRZNs/fjVZYTixbbez3ie6n+YBCeyFi0u/RbgMQZGkX8altzEODTBgi8G95lUJz3qOhdd
2W9MFCQLagYuEp7/YXD1LwmT7u+CU9GGBKHhf/5UF95Rqb0NJ9YEo5FvDezRB+pl45lkYJUrfAON
SBzrWyLzZl+kmFkZGHtLS/ZGaQmVH8gmQLssO9OzAWFmnaiZz92y1BPGIr0OkMtm6nkH21OCpQqR
OqQ7/QMuOIICKHCMInNlM2DAhbJ9rQo4niTRMMUZ1XN0pb0iMnTihnGxmgoWj/rj+/i3/eQxgMIB
/TvMbrhhC3rrrW5tKwluWulEaNlgNQmjwhbF2KjhjFFfpttWGDN0+UFZudw6sZqfLa04S3mGH79w
3AnEWH3WqaRpJ1K9mmtGO+yNkRDlKXkVRd6cYxd2xThYc6R5Y/283oqz/H4fHbz1f7ZEf77HWHJS
BmhsbVOKiPvLb3GFLsllIwPwpJSfubsWf5zh84/NpxkwCbif9mt8Ixkc6kFq/AbA8EJV/Mryup1R
nluMV7WXLjYBnYPDVsG7Qbb8tCHH2BmImiuuJ/fWtUDN4oSxB7wcLkW3H11STC0zGFGh4gSdACFy
+hBxjTE/20aEvMgwMvdDfa0qFmqf7emwoTvjLlPXIFN4kXQxNhI1XbKu0Tki+ah5hwKhmNUbNJBL
2Ie9cebhxv1VQvzTzQz/b6XQKKxoISpGx78Mfn7Hf0fdLjqldg/6iblzlUp0z8d8UHlQEyiYWHAR
4pVZuezlVgQJm3fNOdgU6dDvRtrQ1w4wXsnTUY50J5v19oeC6NKVyf/ZoRAEstLmsxkGFIKVsuwv
wzA5pqA2RZ0HJHeI12welcs7UcupTkJkEFzaADO+5BOEbgGLbLbxneu+BtnrAwiFYKyUPDUnq9DO
oxpgZi+IF3g9jy9pm60Vr68lv9f0k598tmIsgfVrAR6vspcgICtCrRFr43+5AMlCrFplZpRnkhVm
vFDtNK52aR7Mw8gGHVsz8za3YJ4DFHZUcqFHVQc5QJINn9daOz1JDzaIvy0WUHpmlFfRD25Fwfij
R20PfPLT+2m7nLB0xQsHcP5E3yZ9R5fOajtUzTUWPn0lDgfC9N+huayYhQr1lXb8pgrgr+L1dtO5
0EjTAML6tx34520kXDaTsgyIPIh/AcpcTD9hCaObh+g2Ac6690PzRmIuMGKXQAldKZyC5DSDh232
pZokdmELjiFppo9zLzIH+O8iFyYL/9fhzSGEXxFmsCIZUBp/o9LJ9XlthP+QorVQc42j8IG9pEWN
QoxelPKqpQDnohBvx2wMEYWiPC9GACC13ziL2xgPTKJimIMKOa86Mo5edi8Pz0VTDf/5ovXth7Xx
6OO98pX6pgCUlycdeIUUWNwa1oy3QhoLWqcBXkHU+/dd8orEZpSZeLGfU0kkyVSXXG5WjgrDtLXE
N9CF65XXPca1fgUPy8wHI93ErObxr1OhxBNYBvSPogOwbMNZyXtMy6axFJp6Ar6DuGBooJyKDSRg
ZWuFJ6mREC5+i/OZZ7qkxJy5LTSVQ6EB+iLopqC+Lb4gqVMbqzCP1WphdTNj3fcM+1YwEXi/cwAb
9KhyjwXHH76IO785rcL0m6igacMh/XOMSSybZifDSV9xL8E8FegXsscMNBPujE932VjvzKjkUZXa
egnGgtJgpDKJs4loXkyKByOXFk/pSjnXVpmuIJ2jy+D5f1vZ7+8VYYyyvxWzUzF5yk/U64WLN+X/
vpgfVNsNDfHh6jOcGD9zHosMDS1ELYRUBWGD+Y0Sb8vzycmYQAffbBX524efaqnJCJwpj0d18GeG
hqPXDJhblUWP0nM8srJMu3Rod3HjCmptuhDHEWYxUwGgjJyAFR4Fmy16QWSqUc3/7VcL4hIDlOq3
3ThAnI7gNnGEx2QFH8nO7C+O8FMcMupFG/d4x1XP3BMQWmhWX2w0zG68Y8o5/SgAaSP7Ozkpq9t3
yqROTN2vw9QJqAOay9M1nNLAbMVcYO0BKfAAfPn+dFPmCHxV2WcOVlaR5i+mqrMZnVp5bLKoRYjx
X7nt3jO08eQAeKAXFVZOMve67VneRQZ0VZLyu++3UzzOzT0CTVCkCxisjVaV/yegmOWP6QCJ4pdo
LHn5ysQ+6KTpFH2RsfWVsVlMOUSRYF1E3AHWoQEsXrcJ4KuoHRZ4jJ52yI48XERVE0pcfxEhPvNJ
e+qJWujh3W6aXZ1p8unKbu9mP8SmjBYjuubtmntttbdA7aK/weWkV9aOb8QgCr7u5IU/s3eRnAN+
78FIeZjS2qOfvTiwwNQs/zyntUR+FC4+vcr9aBv1hZVnDB9Gs9l9gBRUmb/EXR6FsrD5MSdxI2tK
uaxfryvsz5kl29C6eFY/ZZpxcySK7Tr6K23jdiHwZaOvZLyu5Hu+aOGa5twkoaa5QsyOaAMFZ2qT
QpzUY7nMALVfXJw9Tjq+4ZfwMuFbxRw7T3enUqYIy+ALc6OVqv51bgs2c9m9CAqdBqnc43yjcAhY
CqGq3sDjP9utz20vvgLeQj46U7AM5MVorT62BhzGkss0pCB1FJGz1c4sf4XfhJp5ROsW+lMe44Gq
EZ5RfmvRiYubWDb0u0ZdwooDTbvex5mbpo7RpuuvH3NoPs7SdiUyH6HsLvb4gU8JHvMV8cat5eb1
KpJkSC6I3osX5JcbTE6EmcxKE63QG1I8ES1RalznzmI4247ysLTGbvlAN0ppUXwuHx7MV2LjFVWu
7hCPhN340KH2gmNMlQY4cJmCKqInBZ9GsFAKMq97kz3PKGxLN3WufO2WjTTD9mt2oYJi/9hxpXmU
sXyQo6bZ6kEL4XAU+oT4ihPbdBhdDRiN3wiwX+cay3CRNonp0J1paRwHFECh2K2sC2LUaI1ej/8t
C8mC+ispILRdsVAn7U2DDpCebKvvnjxwwHHgLehtsvDM7AbbrcYWSgyc5t6/w8Bf5SZPK8R+VBSB
ReRRfLUT+XzSJtgKSg5B/0hdZmMnSjsJoUIXuReXfEpzdXVA6joRweGEeqaMxxnA8EL6ybIZVYWh
yUsxtNr1X/0TCbBbTpIIT4Ar9K+WTmp/jnTuk0TfdGxTp2/1NR1Nvw+DWzYnCi2e7TSvMySQLmTk
JcLc6DQyhQy20Avco4yOi7X84aNt/ZR+pwyAQqVGjv8Q9Q9fcgXVl4qyrpSslHYUHjeQ5zZ90L65
Obq1IrtPRr3du1DpRadf8A7Vg6UE1FOENE4l2thH9U/B5xuAEtxj+gVtPHL4bC25BVyI77gQL9gS
Ohha+OuNzOCRs7C0f2rbd0Yge/3L1VsZua3lbImBQ9DVPARALSs7zUI5S+cqf9vKz2u5922MZpyl
xClx9ByNIoqJccNg5+TM9QO750t2gkPCXUK6Z+7nlay1NqWKK71rDrVwHEGlAQg/Fq0eJzZOKywz
UPlGhjHy0jopdW8918PVjUM+Jdt6TPcGEydqYjwY4ZZXfo1EYoVwQ+enBvfDSJQLZHCkgYvyixQt
71MCcWhQkveJ0whGfUgdx5hIDX0mF6KtpGEchUxzbBU7oLRnwVblWL1Iy34Fefp3Gncf7P5/o3z/
2x1piit9rZfhGfdMX71yWdt8JZk4hDYVb5nhkoqx9+/huhGsP+qi1VOWxbgIMGa6tCbSZTlwKflh
OD1TCK14PoJoXOrpSXHXTh90QxsXYT4fBdRmhBTuukaml8NG1nQ1ZsgMRtCWekIDNKG+3BfKafbI
eRQJjHBnP5S+P04V0r6GgTqsuH6UohBAuKU+7UBanhpE+kT4CsuYsl5Gx4CSICZy6dfxV+1KKxTd
1Ii/LlIdkAL0vlpEL6MYv2mheggvgZBUZeAzR70b1g0/bD5E2XSknxwCuEdnM8dcyfy5t2X+XpwH
CKUzqorMB2FGP/zURIAoPvE9l+tfOYfZ5YLgtuYgu8kk6VmShm7UDICgk4U+KYLCOfyt2jMrP0xo
CuTHqOWjXbxUO21F60mz3UHoU3E/3Q5FjeAuWpGg/e7NrSkHtICtjSZ1OHSGLXdRBx2X0hOtDSAe
E1KHw5jIO1jLNSIxKgETFFr8H3z/TnlwBgRcxtGtC4nrTSOqQTjCE7SjdzBiPoYpb3x8TmU3Dn9T
lFRQ3dpMfIRsbpjoyNocJPuNvHqIny7kQTT1n1FycKCVIG8Gi2qhkvv9ENSS89hEZLr8M51kGrVw
F4Fu1ywA3pSPZF0e6R8rr6quAaAEmxbJvoFEnXug1Uyu7yvQFYazGlEMxt/nbOuzd65ejonBes4U
rTIsxmNQidzSny/u2e7lTli6ooG0KpiX/Rjo5Hy6d+J70WRmV6TqlkDQjn+N7bOaRGbk/HI+lq9z
ji2Z/euM/fUmpY484rQkdTTcQlioSmYm1mHCjjpesaoHWrIZ557vz7rZBNWuMBQMBObYgR+CX7no
sp3iEmsCNX5dsq7JooA6nyD+BX4bLqOFGCvbGgl4tIPFjSpWe8vwaCnb0WbuIQ61wurLrTiwL3wX
GTpKgL0/Awfymz1VHtysQ9aU19+Oezdueia80Db8Bm2/DZqp+mEiJSaQECwiRqiZMcjuaeF1dyIb
3tuX1BNOuaAtQi7gArTrzb8r0Q5Jtw+Do5zM4Gnc1X85GjFbD9aMoMA2OlKEl6byVRhhDkaT04ul
9Az6kctvqRO7IMUS/h9hmZDF+KJHDUjKYXBaGfhj3a4AGIxDnmETcxB2QD1N4KldGsIbMFKKc+Yk
RaGbklMJ5cqeWHu84/90pnuHfLBCKC9SdFvzZCqS3Y9UDEGXIn5tZF7AsjIG8hbIK79WJ5RPdUKe
4RMP+uWpt23R9yZqHVFCEWGYItrU5aU/rtDZ7CTanQ8ftTUA+IIxr7krIXJUc3ZkhHve8nPz0yWb
a3n8miZBtCQCMF0I9MrQD4ICTaUV9jLX4uzqIIb4jF2Z1C6BAz1fHicWebR0QbgaQbA/G8WoN22T
vjc+QarBfH1lopY1apf2ylpuVU0wIzpEiP+9PJOheCyuiRrF4XofaN8dVd7qIk48HwAQxJG5+Lia
G8xw3CQGeJUcfgJoXxu30CfzTh9px6WlTWx8SdYRsdKmWc7WCybh7WAzTYtOQ10Yrwry9JbA6zOp
9pk9KRY5H38uD2+sYzn1PMhK6kSyP2eqC59h1tCzegIngDh3iNdSKuyfB8Vr20yRS3Uy6XzoYuAw
5PrSEIUo15vmZZW24U7N8OHyWX4uIrnVRpFXhwoTjB7Dg5hdl9O/wSsscQtO7lEE10P7B80eyElY
a0ahJ1pHm1cGVybrpSA7aeitrX5+mJrd5/RJDFRENRSIo/9HIMEY1g9RSv/8QcU2bXeEgZbhqqbx
HSpwhibGQVmVXk44Owf0F5TBQZ/NX43pMPIWwjIqkOTxpVY5VHBhZP9qW67FqSF4zBOjhD4Nsakn
o54QEHLMGpMEhkboMdalalVVJJDnOOftFua8msbw3yteYaWU36l3cE9NkdxQ+nODwDAhJwd30Dgw
T+hSnMKXUgQHW5LE+9mqylDT85KsQO/d7iehYcxGuc8Am7vqlztQxwulnNYX9C9CpvMlw6Gvp2/N
k3czX4I6E6Dr8oTmo04qvhndLO19w1zxn3BYhBVqVDtkMfnV2ilZ0lN00ieZKx4pxzOLiy7G2bIG
4DUzMDlSGu9/+KqIX74P4mrgqo1HDFTp/7/1Ple6rkUhhOzOLZ9FLsJ2KuP65CCiUwRz6T+gMujb
/Mz0pgKsBLg5nkE3eeiG16mN51tuyauiqGCoNF9GTPwHGElWziIyKJcev/Vw3KmijgLp9iePiPDU
nl4492YSC+qWBj1WjApoSLRYgvoASU0PPyU8HJHuzZKG0pL7+ShqZXufEr5gbPNxZ//w1TjMfnG5
4F6ZzUxMOP+4MMifjM+PrftGbSBPNpfDbmN5UkWP4MAFo+dcg1V4sXXxqbLFbQ3TdFwfG1f/eK4P
hyPsRx3A/nB8aNY3ZkCtJQ5SRUtkUeJ19oDZpSNqu2uDf8YDxQS2zqtbUPhUeW4yPXVQwM1x4gg6
MwX76yukiyDzYTNUjKu5FqeMTjzMHquEKqI5jl442G95Edwq0wsnXiZJDk0ozhsIifY8JYEE5yEU
aVHqB5VtaJN1a/YXVyr3c9wtvMviFPsn8+mNM4DB5UDjb7Lr6p7nachT/8398X3ZQPN2ka3NTXb2
exDTGgQpUt79jBfJdmEr509Qd39QTQAlKn1YXV/F2mQ5Dpo1DE7ix/uYzhgWF6fRyZtnEwUWnKKz
UjUSOyB35p6DheqW27PW0SZbdyCoNg31zhWK5m2Bc7weyBKN05mudRjGShPRQPpkAywRCYnH28n9
0/i/7SXmZ3FhiuWHO/yfjyJ/BloJOTkyQAvnOlcg3vH1EmVYstHg9RIb+8DBLMPmj1H/etlVl1P9
ayrRjaP+KG+8bQKySOodiIpo7bY6q7GIYyW1xBAI1MKzea3jJWgg64UbcHM5cOpiYi4ZhH/XiWiu
BwnT0QdZVg6gYRLULz5piEQnHjpbIVbJdu1EWC052DIo0jykiFhSqV+LGRnSQqKZ1WmvasL4u+IW
B2esKqOiJV93CVdhy1q/HU6Q8m85XEpbn1DnQWKSfyFq3VMV8dYYq9a0FJrYuBUKQWCPaIHf+xis
0C/ohBW7WQRczdWfN6KLxvoXhqMwf80DFnukB5/ntJjP0P1zoMaDM+Ei8Yc8q5xYWNOm4nuW5GbS
WlUzSI2jYXII2tPlCtTUy7Sg/4in72urUSYnolhMq39Fn3nO5tNZjGJfApugNT9MQx2dtDBsFIqs
etPssPLBNYpw040QvmIjvya03yoIE9xFPjs9ERh0e7dkJPsMM9eGQtcCtn6DKqJ/Mja7HJBWkmSI
SOmoQBhXHUx+DoytIIs0rFZ3455RasErZ0cpP5aFmC7JZCRDevDgce/6McQz1GafB3w3HDbyk9xj
HLtlUhYvLkOFOKs8lnHwe04vSyJPO0R55Z/pAiGeJaggR3OPR1szcllPfP7joOXPd4eIMfiR4+K/
HNvz2Htu2vdqvfcP7Gm9lZg+Om/LIEdHjhcWwjAlEA05pXa1or4eqooOe19rAR4NQYneC+C/ZGq0
Ijrkc/hXqXI21VFihaXcFN38EQJ7FRcdL7wv8MSq0vzhEi2KGFhVBldAtPIS62IbLDB+cDmjZMoE
WiXf6230LowWBvlTH+De7BQGrzsVEJJGfyLSVwdAqBpSiTzQb7uMLjLpgL/UJBjNcbUuJ+7d8sGo
QrLB9+9BjRQJ79FJSy/WEQUqsedNl9qfqBqeZwbLxgrYSJg1D/CkF4rJjYuUi8TMHkj3h0E7xHZU
ExPjlWk+ZWbRKI/ZQaJswXCCZGR2X4HMVcssH7zHVNM9XZv0vNggjdlFvOotYwhISW+kPSl6zoqq
kkHDJsM18lbZvjyaO6t2NRO8DMLCZ5uvcMbRFuDA0iVG6d7h5oqmBdsVidG+kD6GiCcx0+sY72u8
wipz8TKOQvxNosJ12c3wlzsSBK3tpkgpVrA0pdKSwTVZvcqeAoE0ZDmDmcs/O11XSvl2TPOtJZae
2Kel4zt7httPkm4VBuw+f5fx74rB06HCNJhCzFlph94zvV822SQuvz86PABfUtCyONXWMMp80T/r
oi+pY9JHJIMaZ4HPUDJZrHyzII6y0WVlA7Vxxcd61CaOtGU4zolyINaHJ+xbz35jXdNrtxDdvIud
XGQUmYWb+WmaIfSnkNIgq6gl3K1vgaj4WMIV+XXd4ye4CMEUU+SHOhekhsveQNknqqvS0golIUSj
15Vx3/XXC1bmrJvBEsi/fMYaw19aZKnrFKt1/EitzHpTlxKOBbYBOBQz8jHgWZ1OTD8ZeYH4BSBg
XCHDkyigut4RK3ns1t53L1Tzgfvyc2U1FUq7jZY+xGBIMJm+G5KRIWp2bebxkqUFv2xUGOHbmKBg
ZXhAiTSaS0W3uds78dL7OU6/Ich0ZyuhQ1bIf2eYnDSRy1iK5XTjF+rYJxrR3vLSqsF5hRDIGiIH
k3+mzW3hIPLVcOyy1LQuqRQUR2pVGEph9kCcH5/bMnlHon6i65z61KwmbkAm2N9C4cqfTS/cyNRX
M5sDn6bJOwb/8pth3c2nPaFWySy8YZ83naxA6O+dJj3s2n7gmJ+a1jr9TlyXzlcT2xcwB+GT28sg
2sDGXL/AVFu0Frg2PPEpGqLrGney/iwaS7iqdicVimntKZy7PU2FKd6Mt3+hI9FuaxkljGC1c/E7
09FcRN0nbVs99mpRSsYh89LpeyrmsVq6Q99zTvofNR+W1wA7ZvCnSmqkIIoJl42wJPCMTsu6gzla
PrUA9nSjSqARo4CWMJSEjpvGpJAE+UKEVk87JCCeLnh+jBiAOYqScE/Cdr70Cm2YTOltMeRjd/AM
Ay5Q0f+4Uxrv3KuL97Z3KnXL5Fx9ZC1jCgMSb9tylUpyCK3PFN5brcd3uQ+JKDHOyHkYlmqd6fa+
H3N6pukRDwkJr0nqBZi+OPzVI/2Kdsp5vVYmhsYZDH33GAoOqVbhFgu2rcyvNd2+aJK9CEC8YX6G
RNrLb6EDMRT3Qi1ImbqEAoaXcZU5tfKF8WfoNfziPbWqMaYeMZJBF6zEe9s3scvzfxP6m1MadAUm
8cAsC7YuDW30bnxSr5dCBlj+piaQ2igCH/4QonxygEDN5WYVA8mUpZUDtEizQg4ATaRWbXjaqGJU
ZWnIN0NKXbxLQeSpjfj1dwQipPVArJ4tTJvctf3q7cb5KAx4+v/vrPbHEVIcYxShE9L6eH6BoSyQ
t6jgL/95KYMUCft0vEc82K/+ImDJKpR+1BUsPfLgheUQSXhqeE4lIhHWiAGilRIMeLn2A81HEC2q
paxrqDz1ewvCVH7s7RL45h/NMO1ktdIIuIwSglDFigPEV5Q2ZR9OuTXcazVDBak+kqaMVSN1Ucac
JqA7gcdhDAmExdpbCjmw5H8EExjeO/Y0Kk7RMY0H45kE/RBzK+FmHlfEn/qFmChEFucRBvOx0ZZT
zeMD5cwYJRUUOjH5T2OSUjog/672NVe5WopmT7PL9RvlTrQ7M5lQvESFQCcxUdV1DXIel2xYW7X4
JQ8Z7hSYwiXjFEq/gaeI3W/21+/V/Z4JVgYV7gs3DyuqSG+K3jDzSbIgfXlmkm2tjDRhM4NoxHTb
6Qr5ZQ4229lLuEy1N3lZM/28ExzDiEakNu0ERu49p7tvuhDlUPR1TA3ZXlj/8/33aLPHzmTDJb5j
J1ww8PTg+L829WOGRo1Dzzqg5b9bDwm3q6pw78VNIWgarCV++w4PyKoSWwAdOwCkqsyJlROXmdxi
25JsQs5rTIW+xAG5g/94QcOivpZy+ssLo5+rJ4kPlMA0P9KHNlHJKhniWU+qadBq6CeGPsnUGqku
GheJOEDNyfxIi2+X8m3sDqw7L56sFYy4j2szs7dOvz6DqCHRWlQ04hUsljbDhLNjqRWV7CcYrweA
SUSgVErj0PAerUgT+FR0mBNPH84sJsOo1W255o4bP9YxEanyAP8ZYe82NsKBcw2yNrDYrRgVsJPq
FemlcI4L8NeEAhwwZdrDwuhvlFANL9dwDObzS9jdJl9YpSEAc6/Oba4vJepJx/PXepaRjJ1IgesH
5tmSKhlcwHj3svvE/QzuKdQwwE7On7B75D80qG4rPbsRsZAZlheiytXNbWO/NskbxkNY8J4r7KYx
vyLEuqRIsR+/lQvkSX6swF7C27Nka1uNlTu7aEB3w7x2M2oea2ZFNlYSLgTBwT0qI5+msGqVvg2p
F1wn/ngds2orbWeY6fdQyVziptyk/0OsM1McFvUl8MrNGpL41UYHbwLb2sIsXo5K2ALWk2wzuYuV
e1q4tQopa5s3CHuhWJa8EClCPiAbei3w06pJgLyP+iTzV4m8kq/ozs2ewn3Frz/+xoiSNW8WkEYv
zuM624cehTf8A9Snhug0zDInz0zxTnyRpZHVvIE3JmFvj1xN5oIEjYS8cdpgPpcj2zX5vzuyacA7
EkWZwSf363vuQJ27cRQo/nt6dAqVNUD3DXtNpoL5fOVI5G+zMTkyuW4ERVyR5p4JcxUzAfG/deKM
9vgpnfRPiljsASCXY/v5rnGnSnYpswb4KPgYV7UrGu0GloyZf2Mb4Mhgrtq1nEPzppddDEeZpEsA
JTBN64deePFGvosDA8qQl0Jwa2Aa3ixu2P44+1EfAzf6yXseHKjNLm1x/xER8RlhlKtQWeTq8QmF
ul101RFw/3ykhDsQZDlLSQ1c82UFODNHeJD7VxKN8FddW4cZXJuv9Uo6DBcLdPP1y1mQfsU0ji8c
2GIf1EUjURLY4eyh6oZTm2QaLQ++YSo1WetUdeAYmvR2cV05hK0TqO/TaiuyAScoXOQKUYbOQGNf
4oUFUJCjqT9MV6/op8TqQeF1/8qaXDGoxIULNmNWeJsBvRn7G8f4zF85y/+cYhwSGoZRr0xQxOjm
5N5+n/CXK2NCR5vtQ3naEU0VmSAcwtoMxadZUEiNs5Ekvo4xrb3LvgGk9WfWUQfDPDyfUHF2T/rs
X2eFBJQaGb8fLrI2Ku7fVlQhGKVmD6YRQ0aLTdyRGoNJlHljnDUfierPFR4dbdlPOA17MQXyyQeD
ewj11f02YePsN/jHgHr5m2wOs+HKSmdq22Js06WNYia3OX+mGMWUCtt9UJoBrnPZx0gxk55c66mJ
DfvxUnRexQSWKNHYarhA43WVv16DBm2KsJbDonFvhnfF9IliVxNZGhcj81mIvbiixNKfaa2draQ1
/6kkadrHw4kxI8H9F9BDyKMCykM2tpYbNDlK8W3sUee4c98TYRyptJ7MGrZTot4D6S3QZFx7GzB1
kDzMR+2YCW3lhu15i2DQ/NsKTHApi3gE8gV0mS9tNgZTEsfqALTyM1m0SWO1z1tqbQYR8VdHOIfu
s0wwHFMv48CdnyuIIeKAT6QprrYsKG+KlOfuC2jx05YNC7xBVZHQ+/eUF4o5+KeBThMwPUYrNx25
p8HRZd2dRePLWONVBPN7DGJuPjg6+rJ2yuqk5XZ8GCbowMMeiFbY8fPFl6P2IR1PcobC0UApeWvL
aduKvf41/1pUoO9anhhp29BewwgdANxBX8EvMJePeD68lf7i6y0Og+gLeCIwEcCSoP6rDWAdE/M6
Q7hEFJWJou7IhCs6PbNPHC0TZtad2lGdnjoXy1STK10l3J8fcVcSVxxvTUy+GYxcVgn3wZ6TvugF
w8xHfAo68mLrtsSccLyD/cbjQRBcI0Sa9gtabhmFslxmN9/edKkSx6sJlnulC1/Sfu0pRPuCpD+I
LDsO0wHj7FFwo/C0iPhBIG+a7GAO11D289Y61auPzAtnpU5LdduqWzEvbrKgYH38t34tewBMuTpb
gOodGzixR4gv5ThQR6a84wmTeu2QKCgq4j1cdCtS6+L46Nbo8V9oUsRWx5iDRtP4d6kLWmBQb80o
UwNO9BqgwYbSmqdUvh+KJo7wTzPC537sLYp9RjGnTEZzrT2EX5EROU4r6tp5eI35CQlNqcsVT8X3
w4RwmnQW6cG6ss/nkIbfErLziugicWxkzawRSXp2tKGKiHHoiDYZ064DSZl+C107LqZT+hYE5EeE
uKjxemEF1b7Pk7jFlf1DTCiGCiAsgvdKtcDA4INBVit17PlKKEUN8H8ye2mStDiaiXMjLCt/0mm5
zypVvJG1j4UfZk8mc0lFH4y1winPC3ms9UaYC4KZRQ9+3YTIKmljo9Sx2+HMq8HHlHYqVE6UPH2y
FFm9VzHWGmt1LyhT0+Oeg7OVsXv/JikJALrBn+3vm9QkusSLZ95m0MZ99BMF0lKfdhMKrowhTXqK
D0gAVi4OtUo0zNJngqVBy9VD0Q8mK1Js8QbKSsv81+xCLQ3ecpU/3nPaEKkf4XxTmFR6GkH0Fs2V
tiAWBZrgTWayo77Jc5JVRMA8NCnwrLskqq4TnANiLlRYNrKOZGjnvnu3mG9ilwP9xg4UCTLMLJqH
6VNTPh53c9ZhYSB93vpQGg+gMVRTM467u8EodG5sOH8VJcgoeuWJHqgLWDJy/q1MLys2Lb6ujXWz
g1lD5rYh4m4jBmOKrdUrCiQG/IMPqFeOqVBCGMQj/KSXhYX9FZXLWkB63ay9uxxdmyfrvQQbI5XS
sAEzW7ol4AW51nCzmfShqzIYmG6Brk4n9V5rIu80PFlwmvOw6m2x9mb1iH77j8bEt/PxWMmVoZBF
iE1fz2lOwqVRprRcpOTG8rczTh5Q06wY/x/DBXTgOZFsZz3K8ZRSVbdUFIVIxq9DMmhYDOa5QIZa
aOY6od1aBeZWD2U5Kha9Y7tW3wGJTzECzqC+f4Yr1U/PbbCf1l4ljQgqdKwvWPnShIcfcd4G7mFv
SrcodQMWOYAnIinURrJDUre+oizR3aM17kipOkk4ImDyTK1rLOFIT+ScEJ+E84flQ55OFxdY7ADY
GmDHAt7rs43WtyDRVTPg7FFeJWiPqFtVfv+DtbQ5Cgr4L8+8bZQ2i7qDfKtqGs6SHjycayQGeEW1
v2kQvfSsUtI4qTDCR3K2mvGesPttnnOCILZUC6quCyEZHnBMqeqAeQqqEKL/Gu9/Uho8e4kwgTaJ
Y/CRs9FMBiMafnrDNO0skK5ElAJFCkKHBMc/VWLuPnLGstZf7uf8RfPpGYRttdYh+cWahCQUjE35
jBwGC1P2MArq4yeOgdWegogFYHfZu+lMDqNEHnupoRqEC9KLLor2kQ4DEcJ8kstjMeSmWlSO2S6L
BasaD3PJAlE1itWOHUIyX1mQsSoRCJPnsrtfFVS1TCt5pdvgQflc+HofvjnpzEMg6m6LYPUNWGIi
sB/Bu68qxTRiyHy+Kiw3ikfYMou3A+BDLb+O0ob2MEUM2HDxzzFOeTpqj1laY3YXl94SovGsetbh
dQ8KNyLOmG9CCvEK413F5469/qR3ddj8uXmdVrGiEpB8SmNmZU6VEuVMCx8WitxKAO9mEt8KUcIY
3nGXmYw2uf4NzRUotIEI4LsXS4PKeBu0N9X4B6WxjqChdPUhctojF/Ay3lesVn16EJtZNeE78I1D
1bKrBJRlXr+66sHGHoIUDPIa32QihcsMTEleVtkFZxhE/1vFb9r/iy+dfMX8Pxxj2Z4Kh8hTSYJ6
4RJw/d8MhjiH4PgBagveeuxqAYRJZ5dGlEOtZTe5FMtaqVYMzFcuQM2/ZPhugpcQOzRBwYKtzmze
0vNRAEC06GLnQ2B02YsSFLq/UIAYX7lfiPrO3UwbnEaRFiDfiyX/gSHsrD0AOkxaxxOJR+JfKeJV
xaJ/RHlZFcs+fAvFauXHv79IOJ5PvvIk9eMCawUq1TO8QezMiUTPfgSV4I9c/yxTBn0WzjCwGHKK
h/6tGzfTwOjyyfsma4SHH55qJ7wlJMIbS+Unp6rwmChi9dln4VmkjsFaBHitmk9LMKviNiXMzq5V
jF1/8xrfpYe8mObraFLYBATzg8D8+gTbsv65VCQxEHo3vyByt8jRhIwENHlmz04fZbz4oa1e9Uke
PRjyBO8wNvUTjk+dFn53C7xeuyxwjXyuYEsDxOBnKO+EmVjYEKBNb0EZ0aGvrGiMv7j1d8+0Jcf6
kQdJN2c3HrhI7UJKNLTR2kjlnUDmLzgG4HPVySFUj9YcytR5GoKiBWwbZ+gWs6dtil4AzK5F4c4O
/eaywc+CIKz1Vf8aBRRqVSnIYu1FENPLfKcQ2vyBP7jKuRAVXcTAH+mZFXxvZuc+96bhuc2e4SjD
uBUAb4FSgmY7Ak4Nq65Vkt8WL7gfIvT3nEhRsRYUODlVUVmzVTaPPYYlwgCW3DdlekrRJeLI97dI
l1fg25nmpDtucpHNPa94HDdjpmZ0HQveqMG0RWhdZHLs3uUXy8DUQL2JPsGRiHBDR01W+IFYTrTL
i1OmZgBcg8owHPIrkSV22tq9fCcEhCDHTy/wf20KAMG+H2imjQjf7vKHAC6s8R0aJGvT8iP397M3
uAW4zDz86wWwyXeRIBl+zPdPyqnsM5BFlvZ93dTfYcv81CezfhSm+8Mqnx6oOe2p633dDARZuN+t
TytwDSrpsVAxKImgLRIi5L+xJyv76lAnANUc7XQsxRtd9aX+tbDlc8bunBUhhTe/Jb5cQXk/jQuH
FAjFHu23suHfcXfNU3hSWJDyKOHudqmbmUPkZ6Se0zXByWmUclbSZohrRl47kU6u2LPkaTsaQatH
R31hjXU/7vPVBoZEgSKUvpgNST99YB4GUCZmeqAh9D00kP+afgwUOV5ucQtD2Gb4rC/SK+3tbgcz
Jog6rGwuCONl7TllO/aYqT30n3UtC1k7b3FPkGkjR4pp7DB17/Umxopfw4VoH+nSs+xu5CxJgkh9
7TyTjuvkjr+nDaKPRvqDLr8LlOoLB+3oacL/BZ81GyRagfrI3y/wcDOtD0rAQll6TJ+gbuI0dIPD
tjGqxMsfh0vsh48Y630PFuTFg/Kzoz2guBhtD+uzbDj03dIrE4GkUGFoPhs1YspfGxn+6fgTtk4m
4ioj1FWhceL5xBmYeEncCL/KTHvy5CwUUbht7vO5JVUJhsaPYNoaISWM14BEJ63E6+wEZhLj8vDf
l2JFHH2VWUatHEWXhWh2+ZWVZvkL8dpcmkygCCrmQEKk2JQ+sS24Wf8ybpw/MYpf7QxGD1NsczjK
xKOUNn+5CGhTVGgAbLydgroLp6jKvcnOMB1+do4HkSQAU0NBNYepsvfT6S5TcugtKS3JhK7oGSnQ
YqYRNjDXpRPRRItkajCTMgGYaL/xODoRf+hQ1kO0UIwJ2kxew1f19knp0u1yaxcyNGJ7mX+JA8qW
RJXmjzshmlZ3e9dVIyN6t3NioTRIWJugVEaKKHUUd/xYQIAMHDTXHZgVKJ7aNx8GvEWRFQmam5Nd
Ry/bX9fgrcas8GE2Sc9295r2B3lbBQ8MlqvZrNkg+nQfmE8S7du4wAlfDeEpyc29e9zPuwFDDZxD
kiDOFTsVTTS1/DVslmIpqqeVXTn8tWdyQi9fZhv6SemH5git92EpolfSOZ/BsGoGxRG9uDGg8j0c
SClGC93qbj/3G6BG0zzafMDP2x5yBlG8qT/Rqd2IfCAWjk7Au6EHyU7z71pwQCF0ttIgk8Xc3V+h
FTel+IZaqIX1rSeTP64/IUZW8mPTvd6NpRahaQRMVN8x6vtia2Mk4LXW6iv3lm81l1snFawvpubC
jvV3fUrLcqBbOnj0zhnt0+wF3AbBrKtpYHG9ESquxpER4TFT/njAiV/MQ3l4RsZNr+oO3ThjZDmi
y1SQg4iaUiRAe+C0vstjY+jU/RiwHvYrALb+tmAcaLAeZXwBsjyTYD9urWG/mFFdZXv1d9feFiWb
92mbI0DGBCgB+QdOFL6m/cBkhJz7jySU2jXvbG3O9y9KCkxnN+MhEO+E7bRHdgr8n4dmOA5e6LNp
gfA6/VhgzkGJ83aNBzjW8EMTh7qm9upvBtSapZjTr6mLtNvj96s9uf6fbJFsajWgJVArF9v406dh
2akjN8CAGjUG7XOQETjafxaCpJK/dACwVC7aCLuWo+VT6Siy00udMn8rI/Lqsxzp+m9ENYz6sl5u
lx/u9t2s1CVYv4i8oKnlQYraVeLiOIz7sz3iiwa7SBiMswWT9DZMjLphZzw6DN2mteAm0Uc3DfFV
ZLs+VT8CpSl8if4Q9wSuVIFFaBxl8StAlqecBaTYms4bPSnLEledNepZlTwXJfpxXNKvLII3bUPA
nr1TjnudYyXwFUyIjgvHMN8z/ppDczevRQznIDGwtGqpURpGUoq6FHwzcZ2OFijVm49AxqI79Avm
8eNEE1GpZtUXHGDQhhV8APzI94lbXedIWoJutdxM6+G1iQyvPdJWFFTFFC53dYp0/6YGwZG5ZHE7
yFWW0UGF4EDSsa9P9HGPaYiaARLqL5EotKXHiGe9LFBqwNGo/PsMzljoAGJcYoGBmbXhDXivuL2E
kMhFxb8//WvZeVy+nmc1VXuYdbawZ4Vr23CMSrblIjzRrg29vev2xB57rHUeWHAufTbX+AfTnd24
gAQBKW5c1STXoH5FIbKibxRuE1pP+FPe84XceRs0gIl6oQl5b95UHL/zUJqrYiUlHmtpiYut3i2u
Ib72EWfKLvWPAmftqwkgYfqnZhbibtNPjdoDVPhbwr684Egn5SGfQQjPtEVnBG7pHpCMpOafWJJn
MWvF7l9CBY0bmjP2FOL/OgoT29bI6yHw7zEejp4u0CO6Ayo1+daprVp9I1GkUWGNgz9MqM0IYIlE
jnehkX4Ok+vyQNcBWIwenHBQz62qX20BHj6M5UZ4xcObWnBARBaSeSg9HLjW+NTiC5OB6Fx+iEOj
GIK7j0isnVvpvY+WF3S2zhcBZ4GHgXXZCF0VuTrhe0u+C3uHoFQS4pLe3bF+8GNiZZcIQwMoZv7T
L5J+zvjJZ0kVahD1Rp+i0GM4ljyD6ei1Jt9bR+kVawwKG78y1Mk0CO6+IemVzLFjnf20pkutWlaX
f4E7SUyZJwOs1rJyMkaLqICdaMdtgAcmm9e7VEKldwyY+pHKL0vCQfM30D1Mxb/1UgBkqCuQ3zsX
sPg1MbppGpphPZTU65Uu4o34hAZMwcKiolgHvVSqlIHlYMEeSE+4J2KxRhpcs011ZaROwKjM9BK0
+96lCGiLTXp+4aTpXyj89XJhpUxsEfED6JZwAZVQxE0OK+YSScdQputLfmqZRDP/FEJm9PUnfFCy
jLzV5PMt121IiXVRY9TBO5VXKNZgWh5PRTfr6XprgXaVRgHbAammWOeR3yiJ+J7nGWfWLEzyOUA1
IgpwmlISgBmhnRfC4MFOmN2ClwY+b/fHmOY/P3qW+xgmbIsvQk3rA2kgUT+9vWdsaY+1cUo0IS48
/djqhk9RKRrY+90eM4h/ICZinhibwHFYWfRMTZmio0GUnDKYIWlqAp39iOSc3FbHbXQ1NtBVupvw
2oggOWZgtR7OFFLEeXgmbFP7plikdl3Aumhjq1woWZzZhJhgzYWilJIZtTvB6dxL9uI9qGjTEjqb
lKNT5xEpJbJK/jlMaCnttnmj46HN3OcJQPzKaCmgZDvmwlSqGYWo58qNXg+c7cZaTZcSXF2+8PCk
bUBjHZNcMLQi/Em9/HoyqozYVnaR0uFKk8hdBBvxFi8TBje/vkVDBomyvXApJLOHOQTMtJLPvPzA
+HZJTfw94fDG/6uGBhPNmqMweX0IWygNG6eep6cZqGyDsovT6NJRNul0lUp2tmtbczDdIvKvx9jq
ffTSy/3FJGRbTMeTcOHDte07nDxsqQOSsteFU1B84LS29IfGyvX9YzhxP6Nhl/35Ulc6gN/Wef6B
CLdWLHNUFWiM68ZEAuXP+3ZJ+K93hcr41NUUXu3xGyPuoKkHNPsfbMMJ6dZeXqzQSX0OaLbYQ/q2
o3N3M6Slgefjs7OLXEbEWO2j6W3BGXYwvBbpVQaQ8lG7NDNu16J0lemyPuoZ4fZiBGTH0DZi+gBX
y0MG+iG6DowzX/dK7qX2cl1f4VjKPG59G+F/L7Rk1Qx0a7XbfmZ0gWNk1MlmzmS542INb1CEJOxl
HcThXONC+1BuhOm+DF9bHsZI1ATS4MElNhu//zgw+kt/WpXz3ZyPDbeW1mnHMWWta08aSyY7HHfx
hFYJwm8mgzcpTsDZaEUAa+YJOo0cKo0bF/uhiyp4FJfKQ2rFPY4MBri+UdmHWSA1tufztAtF+X0b
feM2LwDzeuqlBN7pvGeFp2A5dzbgZ5sNe7laBAmG8IJcWS4ESl6JpJ0wgn5/phxAmE4v+WDc6xWR
IvXjcqWpY/rKVqabgjz4xN0LcQRb1zbiJT0HWxux9hwg0jT+PaYIfCDnXLHNr/csogYRbgOUNvCq
jg1B14aB5mWeJBp+upU6MqTR1mcOxw/tgDrt13BQW1D4O9DWrhf04qqKd4Ft7LxcL+6GBTBsyiu7
TQIQYQLUELOOd+8xhQ61TKTFV/RZh5vZSJZX3UCkhkjBzUurFMyzfKrSfaXFsv4fxymnq8SZXA4m
0H0KFmA10Fs1Kd0oLCWBruKtRs3GGOvyAmQTlIJ5ag3OcTTK6K6VsLg3g9z2lIlplN7VzW9EoD3F
IhU+Qq1LJzEpWDkAGJSKM4u5ZaMufKAzAKZNFZzk8XwHxlmcW2W5Pqj5R6HCxj5wpywrUikuI+tJ
SlJUMVdS5da242NyBuShndTgIACI1M1n6iAxF6hsa2kloYxXrNYd/6EYnwXk5njIMa54fwwkiWhC
z7SFTXzGmQ8Ec+8yJafALJYuaT8kX5FPzfUb6/C8j0LNkJD4rb599zYHS28N2ZyMzPYeZ7t/UlTi
f2QMtvC+rAsot7Qn3VsIfW6GunYPIOccj8+euoz7P08XKI/ICIy8Autsi2YX1s3pknCLhCJjEQY9
STZmvAqI1QKWFCWHmriWWdqeya1MoFlpBrb7BMqiuG/vaL72IvZ5Dmw6bLEuNBU34QWEwEp27EDM
pn6EIZthjW4De760WIM7lhzP0IiwTcTzVx/25G77fb+q+mQ/xj7TTWO15863zr3kCQdogqlxhtR3
ckYGfEFKPSwdr5jP60Kez0/o2CPNbmyNsMU6IQ18sTPeVHnxIBKfHh++3+4rCkYOtKoDpavNFGVg
bUZJNyeV4Fkw9R11oD8vulTWgW58InzrHLoeIjOH1aREwwB4/g1EO0WpLiEZP2BQPqMcwSvqUHL+
ndpljkg5acgpgZVX2AQhjvgCUlGY1Yxk5bNF0g9QgOxKO6CmELfx2axfpSq8prELD8ht71RAONEN
N9Ib+aSnRd1p3ZNQlnr3xSNmZeeM6aZeXjQXRud2FgAlXQ38LrJ4gd7ciQgQmYl2DeOA1aqx7E8B
SykqmzfChCVWVn/uOQAHAog19o1g/E6LZ+5sXPSvKdRAnMl5g+K+wUFWUus3BHGSHsbKEO6kOlsS
qV/sbKcopG6eMureRnHFIjRhEAJ4Hx/gy8R8dtWLmWiY9qy2RYnvEIFdZKrsHpTHZDpeqzF5D6Gh
rtaJ/APtHgCvdFKwfX4gZzM8Y0q29GuYLcuq+XUgDLNaxSu104SbBOWbRqmbAHLQ2DE90uA7AqVx
J2xMYXhn3ykH9yuapbKJRJBk+eY4aWwPiZw9r+1PqqAYV5Iiv0HylzQm3ZFAelMMsqGuN/z6Oc5H
RMT2qRadOngCthPpKyXq+QZBXiHM9cqLso/TNJPsKDQ+xOe7B5W+L20UGfJmgEhk1Piz1IrjurO/
UdduotWS6PLWtKk/r4TCXpFQQEj0dra7CPdZuJeIkoyT+wkAMuLMhwTSGU8uk1ZehsBCwFYU9gRb
zLFO/auslgt+0YMUkSh0bj2c8m0GeG5hiP1jDw7ahhuSI13PgW6bOfswNRgnbx76qA4NAsxFxdq/
s0EO+Ud2IycMiSkMej0nUKJ+phuXh3/c2+f0F77Q/a33p56AMPpGcqlb1fsGvPpyZiHlPQk2vCde
EhdfyGQyDZbzz2shO9KBmD2lMsXbeGb2DV8+MpT9SglYIkcG/QPDvAZLLqTxdl0JjejtIt/rhopI
NvZvhYpJvJOTVpZ+OV6GWCInZIk/2jkMelDHwCOsrDtJXl0nK9MtCCa2Nz+JLjIgNMgdKvABLil0
caydULh66A/2aAcEVr3V+LahWLFGM6j+KXem+WMk6fKiTeVHUcc9MFLOQVX/eZLjxq/0CoCcZnvT
Pmm/kUEQ4o6MQMx3p8L5EEjSoGXtT9PPHuqv3Y1QytQOP8VIR2OHPgLNXPh3L0DwuOFNEjcmSRfb
tF1X90mVZQHSoS0DU03BfBpcgrn/kF6u7fsGC1P/TXl3U74odi/6gLj1JT0Dp2JP2CPdM0m7Qm1r
IS7CyShQX32yzDNSc5fCNK3IALfSbJWNOiCE9xGmRX0uoDjgg1MxoCbnmhbbWj93bsd2+nrlMNFw
P6AxOIdzk3oDqqc2aDL1/o7BcPUxTm0axsPyRS+XTgNn7tuQJHF0QWAVkyefh5Sait2pJarTRcKm
TGJ0cR7Rx3AOc2ZxT1RarLoqR8zK5pKg6JLYwxEU79ZCANnXQQyxrP9xvWf6OZ6hui7eRtvGd+Jl
w91eNMGXXzpYvijR3gKc16u+M1O9YdzVNaTjqI/72Lx8sLNsn9HxGyOmBj1dlwWxzRrqO9b/jV7U
bHh1A+dg6BWHYsbzGaTMlIfKJNZYPY0nrPI/L4Z2gjgERzspBqIegaUCpLaAJtMntT56qPzHiOq8
4DTlAxhwntL2YKKK0JG8fG02Bl8BGHshQ3ilnSfjA+bc6aArCIgF78HRxg+efxRsend1QOWI8QhK
qo0TyS4Z/Twl7JO8K3e9RmckmT5qM/DMg1fok5mzS+0K2O1jEALi452IDpBZv9XWnaRVmBIxKvvv
vQuhmpZps90345dv3+LVe2qkOmOYxEcTKhqQPmhVllMHfrLcHn3nrzQw8TkSeb6C8AemK/peAzUe
0oWpxMICc13KybRC6r6mEc5IqAGcXh0qswBxxiZHV5ZLlFJzl6MepQK677gdZKvjbf5XZJKleehl
gaLCjelTPwaUk8ASs0QgauQ2INwAX8Cumte0++dmG6wRQXfcMoWvGDfgk/+FKXX+sPGOyBLZLWoP
b8FBH5S9jnMtpFwfSqne+Szatt94fBvsuSMEYmYyzdvkBuWYAfBmQomE8y3oYV5XNF0FvJksyMmR
FWgDK9ewFzWMIKf71GgRR/WY6lrJtis/mFxxsImpZRJ4cT2hj/BfLvYxd95UcmEZYJbNWMe71sr6
7k4DODVA30uWIyvxjtN1LIC6V9oW+1fvnzhwWV7jmGgegwfWU9X710ovZ3VwKxfSdQiCJsf0bHvC
tFG/AKdx4PCRPYqbvmCth3CtC79VHEVD7JWjRKgzCzY5e81q8n8FdklfiWw0g2W7vePFEQrNlNW7
BXpeA1511M7X6a/vsFvLtzbc8jEB+98iqreHDz0udZJitxk4EPWpq8XFbAxQ++yv+vc2PA3szNj3
pUMa9RvrPgEDyutByzdxz+KVSprCzhWGxHL0xHdKLrXhrvbWhspaWpxVnPAvyIa9z0RpBp8MLvOB
7gr/V4Q1TU9/noKqyPE5CVSYaZGuHaxShACaHCJLpbhYfLqvNkvj4TeMFlNjlQI24Fm4dHumT0O3
y57jKC/rPneW2Z7PS5wfd1Nr2t6TPkaUtzeFemC3qrPpuxpnScrm1olLrWz9oDegAZbJ5Anu77RR
clRXE+zx1cTt4o+3b7EO5YZoPnfWhl9DNcvWiryiqh05g7FeWw0PfCL/95h4JdVM1sqEoZ6TcD2i
yJD9LKBxoHh5a1bGv8KoQ4ctVTrpVb0QAhKWaXkt3prqI0S6OicqtWpPJVytTn48w9S7bEvqOIYV
OtRRX9wywmbzTql7bWklw2eFC9GbARsduYWmpUz2upNDV71D3YfiAYa1cdbzzIGYfix5YA5bHB72
VChy7DtI7vY8Den7ptNHqbqdYIKiRT+NjmkWi089ZXj3uGUtX0rBuGsJvTs7IHMEOvkEIu1xJA+M
jxHi2MKDXgK7ObPzzkStq15GOjD9wvUUHEiXVdcwtmedzOvoWpOq+ygBxnVecfvE5sO2ur1PJvOK
b8Nbjd1zg3xTicBPHMeCPWtJOpLdOFnFY3+7osSvUw5NYXZ+Fai2JHVuKm3js3aLKCzIdKO+Nk3f
k9roEv8diowSLJgNQCmwf/h+gL/yonsH+aLBfHCMZEwGlDlaR1ogxhvs8+4g56cnbR8hncY/7cIN
F6HPEghK7O2rqDh+cW/m6N5GSAXJI2XXJ5YbIHYduGmaaJ/Kj4Z2bOELaamXq5wF//bZskkzzXG8
RfgTW+DyHA6tnQFKGA8eyA2EZibH6+OWh7RAgvDTgg3zizSrdqeiziJwwA151KZOA9ZHdp2M9cW/
cd4PgmNjf0UrtZqlbLzgxq/7MkiQW1DbRbJcTCAFkRkir89CBdU+mWwtKEYugn8pvVGeDltgyyvf
NpOt6O1EhbKP6fS7WzIbqeAXK5pSxBivheUEYqgvehQ5aQGp2sqagCIb9TClci35IoNdVI2kNwBW
LpVcV5x8oFwhdOssFkw9anjYxRlR1yUKoa8wAr4RV3PHmzw40Mrvtfou53/sf2a3I4oMwecfxzdr
oTAJOS8ilkQwLIp1oMzbpqliTieX32kBRmkwUf36G1BGmzxVAXyfyjNJ1tneCcIKahovim4fIZNJ
xlEYlEHnxRdVkkI8Mpq48sz2J3z81kXr9Zv1Pbmu2gHGFZd6HzYN0XTqLFSzWz6LQwR9EXOIyova
X4hTC8g+zwj39vDX0rETvx1kuZ2uwnlkbixzOdqdMT4cK01MZ7pub4RWTn3u3rrb5B7j+xvLeS4k
wMes5RPa1uEk0QX2qbjvGfrrgnKQ6r5kEOX1v8ychIkAnRauOvRoF6MKkQZkUTz+PBbb9N/Nr2w5
vpo6Kcw5JYPu/QI2gq6Hk66HHA1+cWKKVZ0jR6Ic3dk1XwyXP3d/ABoBiTaSJk8einTOJrclybcI
z6LBZFebGoHPLN7Pp4xGEqAwI9SK9G9GwSPl74hH4EDJr/xWNsyknVrs8L1PsZuootLJt6NdGAj4
+Ey+VGoIz2evqwhBK30Jh5qeg2xb3o7frjYZ+o2wooQrN9WfQSBrYOGsKH26hXmamEyAdbOWV8zx
te8lKUtiyCcnx2IcrasY+C4nM4s2+OzNQp/hNCadwGbSTd509OdZBnAp7U/ORNgnT9CUpjdA0+XJ
4y2i8S6vGbQ7SKhF161yhDyImd0kAB8XoZDZdSQnXCQoC95YIRMv8RvuFEiYF/nl/nQ9K8udUE8k
F0/0GDr4RAV0ysdaEJ4sIQiRbFZLCiqZcm7nhMLqygLXqTXyIZwSKmQDJRiZKFlBvJ/vJWMbUOYO
mt5/di3Z2OUe81g6q5YLz8fcNEHdcachEIMZ2ri3JwuCjdoorjP/ktjaS+xrDFclPVpNYcd14g5f
w7sD0GYMSh5Secspun1drhPd0agAADePK3m3y0FOINmGFoBTaXt/SdiIhJnm8yf5pvGvKJ7qpjr6
4lM47+jG+xjNY4REp//M0emnOIwX/KtIyVQ/ErkAuC8/VpsCD8pix4zEsHRpEAeGNEzzAJSBn4Hl
EwlAJypqd8tsxm+bjCgd8Lx7GSE9qkyDY6pcUHGt3MRBy5Z859FJmTR4ayynn+cNSkVjiY4WJgXS
9MZithaOPZSs/eHMVjiXOeBV29C8zfpJB/z3kWMz88BAeMqHL9dntd1Xd7lFI7iPFA6pH/XGWQGN
1/UYwvoyNABo9tHu4/B/9TcarY/UCrkfAmesoJ9d10gpnCq6GCaBRrXRp1ZxoMug0GwwjPI33qL0
P7d7/utg91LEviU1J9PauMBON1KP1/pOCMXGEZL+CxLOGR5O5xWTPU98nsYIw0QPQSjw189aDNyb
Fm4Idt5NElSRYc5rn9dY79qo1aftpabG5kXoKZf8k25rE+DNU9pIV1QEqBJwFZHIbtEKVdkbTpry
YJK6RdNcBIBVj1wy/odCZ8LEVjHU5hgKKgl6KJu8pJ5Ew2LRsgiWiM4Y+GnOOLSWYwPmJ82FGAK7
ARuhtWjLon1GclTd6rsI6wQ9szqk4LJ2e5i2EWTZJMumrfXJz3KcFvr9i6zXqpytTiRwhbdGjeyk
bfx52CuPwDqy8Q+xfOgj81jMEpbKYnb0ZWCQuxPK648r1xkXBfXcOAgOM0c9HeekHtnO63nwY0k0
gIfbzq/rqJ3VBcGA52jAYhyLr0ZnvEj4HfF3hifVpUDIeydSrqXZ9a+yhvdJb0ti8cMo+ZL/utl+
t/eq40aI9rsnCtY3svIOsNArQABTZTiKE/vj63G0jyYkFKtiITqQldrReitxfBsry7KETJbsflMm
pCKBxzwEpbhQku1R/Dy5XIVZ/L0+HxogNIi3gHxxMdL3plFiEhpMypAiLzsSyK8tzh6FfgMVXMS2
GWe4j9KaQoOz1To7HpnmjZjaT7c/ngOy8Yw/T29sw6WKbDOuzFy7WsTYx6Gtk/75P9/KX5GL+14s
lmUuylTJ1HKIDyXbEeNs4YDL/MDYzSL5Bga9II+aukCN0GvxU9JP4TlrGLuxnvLOnFdTB73ULKPg
1x1PUULJA9hQmIcECBr2/Es7lu75Xbhx8xr7dkmShmvQPzk/2Bxna5TTdpDLTDkXLVnBTgW0XBPl
mdi66eRWBA1kshgI11iF/YwkSEmUqS9+oNDdGd9nR6W3Lj+fIlyVWXYIW42D9ofAZ4hrDvjoVsUU
TwG1dXI0AXiR3dhayHtRc83VxJw+LOtNqWvazWKqfhXJ/lEDSabumcWE1cu5bd0Y+kp4ErosRKvK
pOcwWGTKYZHzwQwKAoWkiTb3pSFIuvrmJlonI65Hh8ZUWEtqp2ZiZhveZbNqnRdFJDbPnfUfsspQ
pQraKjSQGRKN6L0WKkqZZxF8IR6W7nzniyL98rRlJlHFjUAZLc3izLUEKN7wWy6aRb3gjZBuu2fA
Tn9iTB6IDmkLqmThwCZAeUYDgBwK8xKkS5tH32+ScdJ+8EsLkENcW3qLFI/mcQwzESf9EmRgLymr
FwNK1sLXYuo1BJK/SIN3gzpjfB63TbkmVZV5MyH1bDb4MPMgxjd+Bnxa736Pe2k0Gal/7foCTx0k
krFCZJrs5QBcj4ZiDj0zFlaco0p/OVqBXJOOZEydY7ySmo28E1feIFg9fTWkvPvZKQw/Kqv2Daqh
O5Hz4biSdXznzC+EQPGEWVZpG9XoLO/7beaxcujiMzGMy58cS11PgfHsT7DgaPNnYeHVl0LoQR48
x4DqL7SliShVLsPyXL/T9ytlaEgUKgKgxLosVQpUndb41cKR6rral0FPoz9U7BOEUYJAqddIv1N4
14CvrhOBVHdmuYbKNwNZJBZkDr/shUBvHPEZupxFhQq96WiMCzdmF9p4o1gypan/YzvVfVIHFK7y
FnIOvDjJWcyCBJ4QtJx0q3kG0rLZQTOaQctUjrP8y2Jx9VVpZpcqyeUZXLyEnEP+EDe1ha0f8p/R
AYzan35u61oksLC9dW11gaXCaZHcyXQqER26hrj+B8ANw3AHcPYHW6QYAWsSlpNGTnwj+Vv31AmP
zjdj/fu/VG0no8120irKmG4zQGJQzVfQa0r8BOQJNiuHWBvW1cVqldhBTaqYfRVs3E/gyGOqJypS
HcKxq73pJ6rbr+HYJ4dnNORAn2fH23f8VjltE9/OSuECsC7MUv/TOFMGAeAlYiSB/jvqdAt1j/tR
Kf0onn2Xpla0unAK/Y5F0CuB82irSo4kyq48930ehN3ulDjQpSlN5b8ABy6hRjl2tWRU2vxZAO9U
f6PPOLO90Qe3jfN5z+MV/bPdxD8iTgVQfaoC1icUKq5+frmWTuDbb84lzn5bNod988slIHpPgbK1
uBEj6MXTvyQhsCmS054bGxZR347agpKuXttDvsOgm4aLUe/O3gdke+1kiHjygbgYdPcX1wj0LUiS
t4donZcEi6QlUs/JUcVW2YET0oMFXdPsqoDd163oL0DKzA1mxWZ0jPBj3p1/DSmoG/+whjQf92cI
R/C/6jmDC0e9UMsIg9fllWLa5vy5udwiP+KMfg2Xm0Gx712pKiOkJWvrgJLZscoqzhFsLSAlcbTg
0gY/yyPJxf0aL0g4b16DxwsUMzwpH8vfTnY/zUYtCoMHnbCIy4lwKx9vYFM7I86ObQV/HpA0mMA2
p8DfCJTX1Daet+2rchTzfz+grFhtEPqMrgkmDddGVfume3FqG7J6RbviqG05u+/2uad4rwBRUCjF
XeXT1Shug3KTn4wbqaYG6WEpJgoA6jlvfcsuXzSwQNUGLqw/LZrsXPYjjSkbIHSGvbxGGBVPCsE2
uS2mIpRW3ZXBYc06ff1KHU+qaIlTlZRlNYB+K+oW0OXYXo8pbzWw/2DybzwFzoguygbjdqPrMvnN
MsO4UYV9VSZjP6rYlQ+NiSqlJbTZgO6WgDP/qPdpXjnF5k8VSPU+7hW/vuTmLuBhxV1nzB8tZifT
7Lxm6p1YLzaO5n7KhoP8mbUFxTpa0kQwSi8AauG3yLfzQFLaBAayrFMCANSn+xq4efTSjDsEZ+NW
pJItn0EVEoNhlSPj3m8Mj/WQo3AOgFWUhS9JEsS60G0ih+81JPuPKxMiVdrDtPu16/6G9NzCD087
ziK66ZbvTkb/vOiubgvDzRPlMahsMTKQTiv0fys+o2lPvm2ChJatwQQUzQv3FBzTONcDslzBbUVU
FJoePaPlPuNeAEnP0jx23SAly2TkJ2TlRbUGD70gdoXSOzCsPVO6tVa0NTEgxJ086dLG01mGmxJ7
87WfI5KjRXUqjSdsaIEjr0+CsoYLzSefKFNJwPpAM4bcmygEsqLGVA+21Tdzy5ihleHcN1mKKJhi
Z5bSEKhleIkHUhvjCP6X25njC2SP/jgNQJBR4F5ITh7G+YSG5h+RQTWJdf5gcGJgbUqH20y8VzTv
nYJwc9xtCHadrR2nBR/v3OIcubEZSUrpBd/GE6o1zO1LZoihdcGuQ98LxZj0eh92thymy82bQA/A
0975YOqmlbDSjDOx59auLnHfogHMadPP74K9oG2Q3Yt6YYIcyIz6ezzRUMUDasQBG9ijJgNm9VxU
Hrw3gFBa3jnnxz3KYf5pw9m5G8S4NhjIXvZmrCKA+PL+E2zuIrdGI9XBXObGM+6aSUFYDiQX1yQr
eJNfT2BUI5il0QAJsedjvO026IB/LrsebnhnKvWQlCGFFpYWMTiHf+V/SGbaYwDfpLmWL+8MZXEi
ZkuA5Hi390NevcvA3W/Io5K6vuX/OPehI39MfJEBuBXf9bZEAmXp4yLMJMJEdAR0QCLfq4LYE1JO
kebnFWb5kyIxNFLaKXOzQ+Z3qy5eUVUS+LYkQphQoRBSK1BtmGwYQPcDGPtO3hxOHCcPaPhzG+07
mMPUD5rcCJ9UuOLkyngHJ/tsEZ6Zmf7GeYhSZj2kjCyy3ofQxxlTRRXVx9dJRvZKqYSVUocBjtjD
tAJKFxu1KRXi0ar2ag3nUOodeuv6FJl2CBiOCxYbafrX6LZ3abYzWrWyLlZ0Bor2HBnnajPUXs6y
sc1neLcs+FygYGtjo6CecWUooihNm0um78rjOttpqgNeUeotQ9cR3pymjsBr23psXEzgH7o0Ze9u
GENgL486xvEs5q15xPZ+ZRIrr20Q3/D8VjqEoesRMwl5b6XLJiagem5YrsiWg5eyJK98UWMlIpxP
UO+fHYJYUeNjIKMphfCRfc8wZrSBnOSOg5a8sDClKaJH15pD5GYMNisuj6DC129nxYB9f5/jVpmY
nOXNFYrgOUe0xx6PUaLrRKOCbATe2+r5q5g3VaJmKJwPJDhVhF1Hv08QfBMOWtOkXLs5dxe77WMy
ZbR9cOpGIfk9aMnqf5M8wCEI/tsWKx6is3myY4twC8PEV0E0VfYI49gKcsEFruim/bFUleZOq3NF
3yzFudc2TNays1J9qWzPDr5GAfz/gOhH+viRvhJUgjmUAU+zMZvE9W0KtZquIgDWyMm6EXcy3Qw2
LhDmsFoxOQaeF3QeSjwC6PIA4mjRVh+UZ74YvnIdi1xLnybCkaiEBym6sTYH3yZv45ewhilv9E8k
Iglec0YwB7IjOZA0p8GbMBZ5f4QVD3lpoOj8GXAZkAEVo1YFjdlssFA3iaGEkQzgXheVNZLvjTAD
mp22VXAEnrqloq/K8tOQmO2fWu6XYHua1OFrF9QwhXJ10d1ZicBji1hUFBw+Ax2YRi+b1hrgvkZ2
+Hr80iKd+AhMF2Yvde+ekZg+7TIStP75bMlTvRQlDyjNt5sIQjxmsr66TrsmTWzIbpXHYzV0tmgG
zk7ibB200DcbDb3TDFG2/ocok0QvKwOtkly1WXnewkB+0+kI6bYYNgVW9q//90Emg4fyCzA0ApDX
MJJN6vYuL5W2NlR4Nca/KrMjSrr3CBEUIiAJAChnanikAOab8TejsO6XQuo/G92hK94hlttDVcml
XoLH3s2pA6rvWYxXhj90NGf5372ep6P7EjuWW8DqZzXYQztYhjVtsLZPuO2q9dqSxCx4tHVjZgXj
cc6jm8gdEvHNZi5/RlU6d0WkrBj2ZRN+Rw2Rk6Iu7aJKlfG/43Vqr1IeYBVvulQiW3IQg8sV5aSb
3KDhdRn+OVcGeP8K5GW/xdTIPNLwra7XTyUfvz0OsBlIgelvJdBCoW12vBN4+SHQ7+t7ezyEZTzT
qxFhK5k1t9OFBXQ021FcxT80SsAjk0M3m6KwP4fSS4VaKvXEU6s/A4UR70kQIurcornoj5WWQK33
K5Q135qm7R1CZ8ar9P3z4hhIPFfz4ZTR3h9woB7fXqjq5jFJmTWrt12Atq0sWCIdac6RVpH7kr3G
Hk9lEM0JN9niEaiVxAxCTc0fDlETbKGIk1jo/37MzhpyWRSEi9D5R4z3ZTZhMNu7zu0JEzC1jSlZ
9YvFxJIBSJAJzQ8ZET1rfMXO/G9j2YULm0HZ8NpZ76ncI6ArH9Y+i8ypR75Mm+r3B264v50BvHBm
rdCFWB9Ynd/lcKu7k0I2weJOUNKRF7IomTMFhjP3uTWf8Gh0aZ61X+ErbSg3VC6zxvXhnyBYrk44
HUZfJYfRceCBBnFiOkqxTfBVLBU2MPeeOqnJ1lS4fHFAxoTnSYdVVT7KAauM8hhKT5DlpWQk16Je
CUwY9kQDxdST2SR2XBD9r1ZMxCIXtrUPdLtVnkoM1SMvZz5TTDNBMH6yxXJE25YpcVSz8GKUBNoO
wVZxuPjk43chm3Og+AOBkS/FkT6Fimxx7OE4JSr/j/9nrNk+E8wqJXz0OaGAMxsSOFmEKA7tui9c
dX++VwXXSaR5BhCS7SItMJX2v5rjWUG8QIFb0da1vGuEzJY0WdiDWRP3xyIOJkSLm+igz6M6yZxe
Z9N7B++MpXortyHIUrEJtsnsjckjhmQyhq97ON1ZkQfYjJo5+s1X8PMDNNl3fpawXAoDYX4zPUMM
hccS2H0cNr1qpSt30Mi7J1E2PejOD2rKgLV66tjp5h8ry+M7e071PvXn22NNR3qknI4LQkw0dilm
oJgb6kZaKcmN+0yLFfpvhelSTpT4olLE6UslDVk617GBjBP03nxEPhtiVX4CBxj675/5OjngU7vA
kMPces5h44EwZnCfqmWnwe+ooI4b73XERMjw0eVHOQsFfKG4qn493MfoMaHQOQZqoZhpr3JWfMKO
Ee8VtpmWCCc4BmFOtccGlzGZz9T7YW/+oQjCKA01hRt3vA28PtntQt7yC/z299knL0hdbwkmtz0p
7EnMWI12mdkqXzpK86LUwzp6b17VF6F7wBbJEXQ/29Mjy98NSOyptzUnrn0QbtlVfyOvkIQd/M/c
xVSZUK6SeONIKGzPkU2TH7IIipo/O/RSvC+ugvpik2qYy/xuRPOsqbBqbNUAXilaJzBEeUWhOYbp
bmIENXhyU24SgFCfVtWWIPzt+OA4Tsd9cUnlKQELmyAty0Zpr6v+eHtV9ocFy7SsNzWY+yJk7gR2
pL5QQy57Y4AeV2srEHH579CCsmuSfzDOP0s0rEkom0zhbXCFpLCMVLg2MBSPA0FyvE3pk7sKfDAl
cDHrKJLw2Imh0TnyOkQtTsmLcUCmsHMYQtA98eWtfrpQNMckn9FA6KIK4LCsAJX5FUm2AJYJpF8o
I0ufGHSrY96N8+1KYurWIqIL7ep+1cobfJAhjSr7lSh8wzQDZptqdU7IGz6JC80rXXVh4HCgcAzw
BBRzIChVEvGyPjwbrtlq5YHwXZcXrpfhWJCAn19i0eVMmYyNsCLwHETH03Y/MorAjfbXVBx7TvPr
YQEPI9Ubx0Zd4f7x0BufCYicaWsxfuikJnio+FkYDQwN/lhnkoB49Zc8YTa6H827jQtfWVlK+DJU
+gsy6ExWLhQ27zKAr6lNIuUCup3LSUskvf32GUuavAst+1h6CvqAYaxUudKvuJBea9v2DbXrYnVl
M40YQqLjMbpi1rdTAacHSoABBuXHSSyvwVpyr9ngculFTrUP3va8GIAJINBqmUc33yXzzcJpD2ZK
AuiqbI6evpL8N04mtgOsq7agdGOeiyRJtUy4q5/td4KvKf4p6S5RJvhAHNqo9+aNsaMhyDpaRbDf
ApgmzJxHXM4JGKmUTXXaf2bNcQpo8B75UI+MCEhHJ7tUzNAaecNLDOiOP9MlY2uw5IxK0txTfC3e
fDSX2lUkhYLNYhNaHzdZXO6sPUK6+dq4/G73AXCL2kLUDF1bM/5Zw7S0dNUzM3gHyM0zW7BdUb6T
bs1LnRYOG6DEEFd2QlDdwDEg5/ZBNO0aVvsyE/AkHA5WWIlmtvOA5y78IPLRudyAntlfcVdYjJ5O
EZEsDT9hFnJRraPQpDJtBw3mf+QHU5IMjeSCtw/qxtp4XHupQIYK6pgXnr9qPRUCgPSWnJtxveFb
nYFXhYlzVcbuEkB5MpQxX98sm1t8ovAvZRqaz1cqnw+yQXgPO3YeTyDBO9uGQhjIG4PJm+Kuh0zd
ictfW5sGyiZHZEMFCqMcwoWJXWVwk20j/roZJJLBNRAuqyCk7GGvqsGWhGX0SLYT9RTdod4U3SxR
Wh7tQg8DDbXBsw5kgnLyCD4x1Y9DjAYYa/CIb3XKgOy7XXniILodcVNAK2OUatQ1CBUsiX/GH277
XIUeHUbko43gdLW92lNqMo8mt0ZkljU4BNBjAie96NDnpH2NWuGWck0oaE6RH3K12Vayv2cXYtqg
n0QrSHayNAoiGXjHPTL6xB9n2123uTbQj5EifxEAyM4bCOaSyv0OIZUILgbPm+XVW/9T4xGOIUnd
MNOYSlhnKGZ84SrT506BIRnHbSUM4D8+lVmc0v7bqniP9cDNvZL8VfglgPGYpkzWOeuSD1fGPUie
eikbpbF0VWEU1l0iZ6JYVqkEs2md8+w0y4tz5x7Y0yNQvsCGAcnrH0doTBFpPgxQYZycidB5xgLw
+6RJ25vaZxfReu6gObIEZ+w25pYcLNv2sbuH0AKg3PIwpcNTfTrjkfmjMWYvQT8Xl3DcAoV3//bV
pOSGu4zanzYeNI4QBoREpQYn8G2+fESRcoAuTG0gePDy99Fs/HsmrNBLH61oTYyX3VCQednNIFzs
qB/WnDW9TNIaXkBUgid3lFSTKHMyOFMwH5IWtyBNMXekp9FXP6tHnZ59T8bDHc+5ASa9N0hDnR6B
Kqujxl8b1QmEZiv02eHKeWH5M+urpAw6+02O2xffHRRBGO3iRZDKCYYLecLSDr0E44VTJC1RoyD+
7EZoU5ThwuU9Cy1NRBEreUjeARp5NFF1+8v4yfc6G6kZhZVNq2eimf8F27gxBLJfxbdnJRYTTO0o
+js/s+afoY32a6r0tfKNe25lU4sQhNm5OnOOxRS1g4UwjjtOexKL45E/YKb6pNPZ3jrf9UlBrcBG
zlQwXFzq9yx4olDdVC6MOIsICx5YWS82HfWMCjaxbavzVafjvpCHnvzoUnuiQa/gncum9L6JjZd4
Dbv4+vMXJzquAtbpsEnIruDaUbbm1E0B5gQ6ccxfnW5Hu5MZZLPd3DzLZFLRRWBljExPCHbVDfvi
ABNa5voYp9+y3SmJam0JnJO7etbjIzIwx1sceqG0Se3LeeWzHl5yR8OcIylUuR6orKe8gXM9Ps+W
ftikk+5bDe3glg60yqAiEygTmlsiumEHzzcUNOlsN5GJTy5fu2NMpq+G1r7WIwD76g6zwJ3wMDf6
ZPJDpF96eFQNRESVNksmVB41TchiKGrjzsMGDVOwJrgjrwSgmEURHXIeCTOOyA3HmVVfzuq3ALUi
ttoJC9t7sGoMm1b3zNKoOJoy3RSX2yF28tJI5yCNv6dl95Ec1hQdksK34y3d/tRHXj9pTxN00oqZ
11UM2VRqShsDoxw3xjUvFdP6ju8WF+xHC+pEsNoshAzRpnBskMAb2W70LteoQ5CS51RgQj6wvxaE
gbC7JN45iqWplva1LB4pYL1Ydl7hG3fQzYP7sUn8QtTbewawpWNUrQDx2oBe1pGujl2ya4a6y72q
wKrqyzbRyNmWEJnOmuiw6MZRaEfHPrjehY46KVVcUZ1fcE75e/a1nCw0lTVTSwuRjDlG5lFx3KuM
Scnqpkx/gAiVP8MpVEwAaLN5puXEaVjiI5jnTX5RqfWHCnqmIbaUxA+7How7LPP9tQhMMflDSerD
aPBXzofUp4R/AK9ARcorZnN03CYaMmj/Of0MYSu1yijdJtB6WQ9WYguhdlZw2ltjYsMinmYhMO3O
NVek8Rew04jk87x/P7BJJ8grL+t0x+pNsd48jQ1EPkEASnSwTdGmXiXEsFFqm0+ThS6y5d+Ra81M
EfeNt9xsRChYABq5/NUFT/Lv8V9gDiq5Ex8bDPQwaUNhRO8ARAg59NuVc6S6GIrBU9N7xuLZRpiD
9RZ6agABeffeDpmudP3rE/2hFoWs0ZyWrvBT2JXhRH2mAmDyD65tIELv4BbR1KSjc0936I326Y0b
rsJyUf8HBOrWqPU1aLb03unX71XlioqDzxYkOkgxmayIXiD9IkJHNA4c/cBCkK8SYgadGluMkoQ2
pm0wi4IJJMV4wBeQorJteZsCfXOFEEy7/OXDI5lO7orozLYI9Z/mOJrUI5Y48N8kfZFZH/yewubV
qARO7qw/XcCIJK8cXVG2CLO+rJ4uj4ASlF7+S7EP5YyaB8YPWiqFvHZr5GuH3ufvJqwK917LCL/j
dUF/qJl54vo/9z0j1ST10z4Orswj5Fnw2MRT/aEnrKgG2x9t9m5Z6dUWJX8HVEdA6FKQPr9xikLH
vkIALfkFc17Dmbh8LETSIGBf9YGtjFVPuU2UXip/gUPDWB8BY1JvUBYTLmyA/b6Yid5KlT8inNwc
H9CHdPA+GmColODT23xrVCHzKdOKcwL3RuDsTCzLWpEB45cpbCk3Yq9Vgoqok1gnMwa1vkGdB+vO
YzvZRxiG8FsFq04i71zxVzIruVBSQpGYgRnWZCMqG8W5QMSuDk2dMd0GWN2PGGH63wCzTNdtP5JP
gYX/OSQjNima8aoM5CMbKvwE9xVNDu8MOcal/qoPbdFI0v9hzokWaftH5VjP9wleZu3d+IUWpuvU
cAZbmxhCDlWRiPoAdJFoRxTueU6i49SSeUbp/gm9PjHpIBoqUJEb8hWwS6vsjyWTTQuEu2vooUri
2eWdeVQFa8KSYYXbJNDp/VeKPJZS9+g8TflbkXC0lShBaDIrSjMVH3g54ELuIyxqQCOoBOeybRbT
EOoMvEirYEuWYJJebrgdB00Fh8TKLdw8y9Cc7AR8SB8aRRgd4X2I9+jjnHSmXONozyi31SJ/c7Em
kqH9qGGa+OkR3xdy0EkvgDjt+KAsxHHkufakoQNFBgGOEN+Q1c8UlWvEWmjqY5EnBGWqYlxnsI2L
y2SWFjmzQi+smb3bAWbdlrPoKQh+BhbbQR1Gl7FyvA/KG1KBJs3sUvK+fo93cYo8XKyJkONDaOA4
vOjEAvjDiwB2ZovzB/eYgRhhsnRIbcB/eYqT6iaxsL2pvy1crn3IkNSwzpUERjAI9+1Py34vBHNG
BcJhHU4btDFlKUTss1axSeZxNHRnmC6p/mLaxMOlE2yFur+fFfG45fwNsZl/Yrm2OWSdbxCoqHOX
1Yh6BwKwLr0l9YAN56mUCndb3FSw4UsEoG9eEFOvthUubymApwIb9DAkn137QpGDvmOhQS8KdUXi
S0b3kW2X/KnmJ39oasoXJCEgQGRhUcKPsRI1paE47sPGMxz7MwE3S3Qh20ukTHAWLEINhcHRAAfg
C/Xkcc1EDJwG9pjLpxe7Eyyp57WAerAhEdSOJXhfRVMAHqaK/nBo4nLNskz0zJ/nX18nJqKnStTH
el8fg1iLSbPZXmjVQlLS7Oc+7I10PVhZvVxCGMlfaEx3X40n+ByLF6+SZI8Ej7AH/VOFZrIVVj9t
MQMAFJB/Zdg3VpLeiOi6H+H7nlfMmPnD6g/VI48s3p/3n/BVxTpqAsfu/+S2DNZjI0aYw14lvAma
8yOr/S31OzdmgFW6gcDY0SN4tANrpXdonM+abaEs9MYCP+JXzOWFGzpfKc0EKPcyFwbIX94Okzt+
D73FKMIa5PqGajJXqRXHUTdyWCv7jLRgoPWMAmBLrTbFRHvbQs+S4asxVO+h4ihApgzi4QldtytC
R/CzGIJbViT8wMNWUj4ZXly6T24mHsiVzRm+Umb41byYML4AUOMWHEFRUpSmJqUh5p9F2b5r7rhs
XyfM0EvaoBqf4Q/8TgsjxrfnnokvjCRwuQaZtUlgBi7oS325OkfgJP69RY69SdwkXGVNCdDe3OF4
7OyYUuPhUHb1vGMQ3ga+qd4ztJSWfryT2K3wo//0W3u6fkG3EFZhBeS8GFcJWYnvca3exfaYiksp
fBJXIkf3Vg6aodBnUHQB5RG5LAywlrvdhOObzeGNbXI7xaew2uGqkrobnpHPAI8wl7PDcyje3zbN
HpRomgV+VH9vrNzi/bzJIPjB4HcJioqeX2b/bwhaLIaRpROCF/yDOEoM2D5IHCFbm1Ih2P4CLyoY
g+mH0TFvNg7ecEnXSYOr+W4V25GB8QZPmzlIr/d/ukmFr+a7olflElimxc930az+389S2XCJ9ZLz
H7egcSlIBWHUTySm5/b3VWkKhkeH3d4YLUBmWN8vp45ruGRVE6DjbPEcQ3n7PqsT1LdjsdiZYkwd
9Lf+rz2+LpsKuA2R8acozSCDhIGLJt8JOpgv4vpRcXjveAWktrXOEBf7os4cwk9X4mdSTcyPxH7Z
eNdIc7UmtaRcVKoeNGqdw1DpWOy9KbkXcc6e9WoSdAPdZ0Iq1fBdUdLY4do2AgE6XS50ewbx3OPJ
ZvHsfOjZX5LkYZ/RdFolQKWQ7ibXqQbIdTuxRtm/6leYldozRzUfx5aIbwUdBpMNZR/4tv8Kg4w+
kzdUSby5K11dYIYjbG8QDD7W9KId22HZGlq6NQZVUfzPyNOXrS+l5ATM27iYVC/fNNkjMLq5J6Yu
a0humsR41LQkbfoGO988kKCGPyHAMCskqoq7xm4gwJDPABgl/OFISDcscDmGxYQnuKXTloQEIqBt
jx8iX+c78Qcqtgv8dP2kV2NI8xckGH7rq6TRyFO3kAKNlngN0/NQLoVz5f5Ejp/ESg0bpF2canWj
e6+o2y+F9iz5hdkzb9BdfXWQGnx3V8I7nWdYdvtZBAXFpgU20oULA4MIFYxUkr/Jpoeq+WWvoQy0
6z+UA3/BRldBHI7fqiL6JaGVXHhoQk4BPNC080pGbfuNS9iVEoA9nW26xdfjVd81Rd3QtsL4Qnjt
q6uPgQZWqbdPbUYorRBzgz1TddkK7P2fuPqmkaJpcahEmnjrImyFiUSJ2GEltycBeu0yd5QRaY+w
Z80IvbTm5tK2Nt9XUYfq3+htzwre5O6qSllutWdZc8llvTgvcG1+7wJyTimsc7bhqAF1np3SkykA
+mumaf9+8XcxSg48eaQxvC62/DrZdiExYOLXUIs3GNfAAJ+6d1Y5GiEXkZgd+bj63MSQcJIipM+2
Q26ACQ2KxhlEWPRJPC8VDPFTKtvVJSTyn16frC3lMLsq/U/JNNCwSv3DUspVepj+kWy+VYhkOFbP
inhZvlFJ+X4pGoioJC6PeBAI7ks+KZwCLpqpA8QYXgupdsaPV4jmN/+SC3RMEB5GyWm5BRgKmUth
40tOjILB3U6Bo/PkbdndMEE4Y7RjdnFNZYPBgPNFfibQExXizdAfdWtuYlqSq7C6PygyVcQIF6Ne
BQHHqqtssStdv5ykxUhzZvb3i0ttjl8a4g/862Fnbp/IKDh+ZHnO2KY3hDTO2nR9FfEWkEbPwQE8
tv9I83fzp1HzaaXOT82dB5rcxHKq/cG16MOuZuML7JfI42gvWs+Ds340YyURuC4WNBtefeJN2en1
geDA9SZO3J6X0/Uwse2dPMa2/qniSalKGIxZ27DZnsLlyBqwwT32WH8Icyc/tKkfxobatEsVhlkZ
pxMzp+xQ9sKrsXXg8yHJYKDkxZIr+XIE41fBn37GXNOiAVVXmzvW/Bq3EXArkmF04YrAZtmXVDSk
N8GLqc8d1WKl4heZUoO/s6SQ5oOB7SNNuyqJ0DxUFH37nxpQpX5MbFm04f1zbucHXtUrK/o/pm4F
7+3/S3ZdNN8vTmHvUOJBroeGvGrGZ+cIijbIHYU8yjR93wOX//i87TlA0hSxJtUlHSRK6qrzgZyW
qCSut8O1k6eWSZkzVdNik3eCMeB5e3UZq+7FuLpHvBW3CAuGF0lzomFRwCArCaD+1h2qaxmLASDK
VZQ5hdl5k14/F+E7dKE09eSspEMza6UjvLwS2raDCTDbAK66ohRdZGjkwzY77pFoCOKB40GbKDX6
146jzsuFcoDAfteNATIqYnSLQPyzmfYxXqvujX53bC2Azzv47/IJ05qf8vURhAPE0BY7uRvmHVcN
ElbRzt4UH3ph/QTbcjfd7nd2SRmQPct6J7evPLQrtQTCR0R9wcV1CUyZeY6dHP8yjzqmVSlnxedb
bcOcsrLoDeM+OpogdqVwDhGjQT9J62uU+jLvAAQbg0JwrPzwskjHmS+QW0HsktoH8BiwQTgKukUk
tWYNjMbBtpJuWjtwKwCE0unc9abcFBdIxHwsUdM3QsYa6gEqkwstLv0pqij4GltlLuieO1dxV9K+
Dzc9kVz29yyxvCuTj3O38MNAMuBqVVFUCAdVvdvwCcE2myoHGi10mbJjfL4yAVLtaLCY/2L0KRkJ
wuGOW07AFdPAFGF+Ukm38R2hjYKwxNQSYG4BqjpRY+aSTsPYoX1UThnpR6bxxPoMn+XNSk6RFfTd
2wxa3DwCfizpiEt8Oj7ueobKkyXMPQPcLdbePjnTmTRxOCkeTiNA+FARi37YQ0tPWrrhEBggrUmT
LAioboJTYYXVmpww3tFRxBkgAH6ao6gzyDn4C1qUunx1T1/zUQmzdcRUCW683MkpXjYGvsd6IqEQ
44EpR5eh9K4KREusEGO5jSIVY9CN9FFEoCAg0+SkqPeA2MiWpL4XNLHhqwCD9Zmea0/k0qYEAAC0
d+1/U8pt0HC3jNt0oEeRoyB4Tk/WUfbdjkGrJP8WCDd1u1UjpdiGiWuEMnuO+Sfw62W0xXmmx3aS
uL2gh4nEvt6bb3l5C69szEpCzdl1O+ijyZheW+58Pb0pgq9+k1USrsQL38DR/4L9tKKQN38mj5/V
hm6zVRU1CwZ4M48KnvsmXfYtw++SWhtIzq8KvjEj5V46JBnB6nzcThUQs75mCtv8gjJNnD4vO43Z
AgrWBzwJHn7cjOdtXv/iyqv6k1PVYMGqRIe8pM3GIHfS8i617fVoDilTD1a8tJ7hp0XHnYwMdOf0
7R1jrhZwmKCtNJnGR8sffpvFOjrhuo2nvwCDxXUVXp8OeAiMXS515gF1kEus+lu4fjrwjft0VcJ4
8oh97norEdKdu9zWBNcdbDX0XFuRkevd7AohqIlzDliYHuuQatJSY6mTj3AKpBwqQCaxahCX3511
YDCOvauFE4st7P4nIb9syjvMf7TJSd5dpOj+sKIFJAkTTIYh4zXJvGOxQtIQ8gZoavdC3FZxYeWZ
mWlM9+OPB4szi0wtd4isvbL5PG1u5+b0QZZ6YvpyU3A957pUZs2/z6rjbtNL53aIvAu+/fdXe2L4
OynjJ9Oy2t+zHyY2XcbrvhdqOLW00L41uh3oOAN6rrhVqSd6Q1Rw6lBVOgSVXYOqtya6ZmSlto1z
5M+OWurZhTPMfvcU2Dh08rb/KcMFrBr7pHGi53FY/r40Lx7CrExZX+xgTJUZCbZ7QKCumPPvUIvN
OEZ4fQm0poN8wntjyKLbhNpLslFIcWMWlvrdrAu6PbZ2pmy6vxod8qaOiVp6Dyhy+Iidua1OBeAx
xblulWEiNb1w4yxs3AgA4YZkHXqJ47TxBnPIYBPxz3d6thVJnkULCDyZZc59iG4R2B2MAOtUmAL/
4hGRRa3WvFm6ceJzTcKOXxEVs17U6MEE4RoytbQfVn4T9e7C3fsgAZaij2E+M8YCVB8bntj8K69W
e/A7W/uw3UUhAXHjK5OtW9L1oH9BXUXiJ87UERojxG+zzC8QyUUrGXQEfIXdySzelJYazFl16ksJ
j7BK0CHSeKhbzPyKC0y+LP2GGmJffcF0fl4bbY7QYPl4V8UV0W6Qq1bQY3WZzHgabuqbP6lptPKU
IO9A4jJ1NCwb1uWY1i/sXrGrcDopXYkBL4eNpDZZVlizZthtpkHXR7M0TMSkIgmoSZWUpXMKANtU
oL+bdULoNA9wi+PPXx7Rb/I67x3krf4xl/KUjsrH3cJmYcYXEUr00MxUf5w8yM4qMg1aXePmeTe+
jB4ax8s7Rt1OwLUzDORyMEi9dheQgzq+9u3yTBBnGQbSSQYndt/hB4Conmx19S/VBWCzblx/tl1s
QLwiQPHvFmr8UkeZzCP6jV2vSjeJRXkhwNzmPM48YSFZlQpj2Y2u17Vfth2RuZljmQlw0M5jfjhu
aW0zQHvEB2XrGAhSy3eQoeNNd/l6VsmUkHwb6sQ2/MsMuA9SO7o4PKXAINgNzO2mAfdHSTyWCc4i
LQU/2111ELr0qzHmF+UG/DVXWJz9zg5gFVi0G+tuOekY3r8nEdyZI0mM0C8Q1OdB1M25kq44todO
tMA5Ns38uOiPg1goiquFsgJDjvTLyyXtXYhrrHzw5kudmmgx+rCiZZ8qCUn8Bh01qEH36u8SxrBV
QwxQkRvVfGRbVeiJzrdrGkXrXiFadgCYrFdWYitBOtBuVSXs0RhzRWSsluGWKhgeMOvaYv+M979q
Vs0YPseuAnZxOAbUGKWD7whCc12RWsbHhxle0tHycjNV53aKDtA6aosF+AkHQqVGjGgzHw/w3j7C
UpADs9DlpJJjRT5AOFwxKWIfy17lN1wLeV1aef2dMPAFX0AeNrR4nIfqrerREoqVIVwUsuX54L3u
Wu+4i5b9f/TYi1RydNw8AJrjOgSimx42/2Wt1q1oB+0m+bzoDfnWDMhhtQsja2TDh3tyMXmAGY1c
Bdt6aTPsnGLSlDKdeUvCSftp67jyw6aIDrpPJlfzME4kaWoGyzhA7s/PJqluubGJ4SnuKL0fwCWB
0v6Hn6nCA9EYmfzp0AL2v6WKvnNFjCEFV5FWT46wp1Q0FWdf/HydE4COvRuyxCYG5P0hSS7AD4DH
0IaAalip3ob66RQMEe1EL00G+kFTLb/LjQVjkBKWDXDkBbj3o8RxjZOXGCmfPCwLk/dusdr5sRha
V3m9CCC17P0IyvEw6v0tupFGXudLEEqk0M00wO6jSqQj/m1aSZBOSdntZcN/yBGh3wdlDsdA1lf3
VstDt52a5fncFHEj7awNpcjOaV2254SxErLGJBdBPtP4pPgtN7xTBS+DFyoy7HOafspZACaW/Lch
sCPfKypvhmmOSpx89eeJKjAzmpAwowBmVGe1qUZX8uiCw2dipksIQ2xseE2zu5dBydMAP+Yl+cYB
kUern6Qb2OqMDiJeOuRAy9EBSC7iW9oFImXAyMojnl2G5ngHhUeX4skGQvjrpvocDlft28ZCCEj/
dQINSKDG6BcJrCvjufuyiheOu1ElnVJg2RzXtdDi3165bD3Nxgcw0Ta087/9iEEBx5zGJLRmshNl
QnXhKW3dtM7etXZn8nGhdE393GFjEa4OJYBwSmhOQQABzMa14F41PzcHmQztDMPB7t+79W3Vo6ic
FHgbOzU3i+AVvcW0r9Oeamaz+juXJ1gFfAwHfufDhQhP3PFeZArMf6X58E+Wk4AMOBcP/W5kSw2N
B/D/7a1zcUhACA+fH3z8wttw4mfA4AivbwpO6YFvJ8vJLOKewSDOxbenfS5ItvRj6Fb/bMZjoj+k
1DTlHBhicfllagnSmc2QKQFY/hbCTHjN0UMtfi9gLZ2yqWOm5cFsS5BnjIXQX9iZJZP2CKKaGoX4
i6EDWxC/LaAo0KzfYqM9kqMHDzhSg2JSgdtYMryOCDnxevaLKWlqIMm7XAGiDiyt7g1Z679Mdy45
Z7bxZxNOl3J4UZ1hyaPprBVJsOngpyTe8IbDOSHmnKN33R6luaLDogjNTI2vSYKVxr9wX2hS8uOz
52ON/cqhAz2EF/bHQAkOu2wUuPXCjxiWKTYfvxFj1+5cPoRBht5EU/9FwJESD0CYxkLcuf4JTaZ6
sr15eNsGHCDlJxPS7AyFyOCA9r+GoNZf5wzgA2aVXU4e5Y9re7opmisLZgPJdwNoWOit9inb0F4k
ViPO9pJYq4QgmJiYLSgQEp47Xetj4fGfMiDyV59qf/Eh6gZupC0V0hAd9kWlfIOmUlMxy6YfByNO
ni4AqAW6U8RUIXwOkEE3/9sOHlwGj11/BN8rRrI2brZ87V+z/dKsHgyf/DeIlt3h2Ur1YhAXmu7r
5tLXmvdZ8iyCmwR4qh1dZBO/BeGeEblqAWVYELGixevgbYxHZzccetDCqsNWd6JCN3Qf5wmEsZR4
vhjtypErF6tdU8ggMDK+MhWtMvTs4/gCRl+fT/ZCyPpFwiAs0Kthf0+YxGZRl59Fuv7215KaF9LE
rf1z9c5ZueCm2pmAEG5sZ+WRmv+vCxkT99BUdMgnIwvXyzoRxj95MgtZBRJ6QtyjbFJSWoc7fmSK
IjkBeium7liBH+fRfFmcTSkDKhYt41tGxu+i2q21ZRfzhYnd6d3vLIHIi9u/mGbHHnQcunjazO9y
LsydqX777xRfsvr615zQXARw71vHWseQ/6a1/QzLQqISES6kapZFTZaRNqAYddBhkAx3keNZeshF
3Q+KysmgkSvfQiKKr96oRuD0iPr4frSmp8d0ZNIDcicXx+PglWHYUS2CK6srEFUMkeMSZuCDEx8b
u9/Z4i04W+VTrUcnCrIZJOyVCxa5wZ16bbKwyvbZoeXYsTzT6efNgqihX2TACYq++4mXGemE1mUJ
tlRj9vST/XpsARQzFDJSfFP4l4KioArZMKoI1qFp16oMOtphUTQZ6aVPRLOLaEGWi9AbHZ+68eHl
rYudDAGscusnzr0NaMd9Me7+xeV18tRPFi2bzDUtnMH8N0aPitrxEJlU6W+SA4nXzJv42iyeP3h7
ch19Jj9YS2/wGDh/NGXbMah8H+p5zu0/yKeUAtpoUSSgR0JNZ/GW2oNcIVB5kjMMNaKmkqyn9AwA
Poj+m2QGlXpnXA0o7Q2Dx7tJFZskUVxOb1ECKZQ7lCGS3+3g6TXx+ehkBaTu+KDJs64f9OF5o+qy
73zRWBBbA/D+q+KGuz6ved2I2Wvvv9hNf9UJkymzMuxQG6dB8ejmGoaI6c1+f217G2NsDg5rIMic
Gq17Xa52g0C6JbGjwAzsDNd7fjZ1oQH5ui9JwelDmr+ARZtY1fxz35ImS1d/lbluBI5rezHZuPIJ
wFaP6RjfX6rFHBFPXY1p7f0RL6YHIUKVN4h9fADLp+MNYgyuBe1KkI3NeKUBrtDrCxz/nhvmBlPD
KiR2Y7WG+PZY5IwYUMr6qfTqixzsshFm0AnHZsGCShUqKFMnfLEuQScGmvhXWXM6gC+Zi0PMCOIZ
AOIDFq1kUyQP0IdZ/5cSE+NLyEnt/QUBtexn/q66k9AgxcPEzS3hJmhUHtMaPraKxqmF427jtUS+
e85/8IE91PBiyH6vL4eraSoReI/h6UJsNXtRmHCaMI3kkgTElG7zDx7kAAdsXp1HZoW7Pz2P2J+O
RtSf4bSrtocNM3Z9e+o8GZm2NiXgNfuyMaFjEab6Nd52RCIBKJkfcKnJ3BxhUcFdm+hRXbWi9LJq
jVcs+kagmXYYwP8YnHzTO5Cw1Jif6Fvij9KIny9wqBbltU2tX4OsaxngDW5hYEOjsai+kGkDLGlM
3+tzTBRvGkHMgpO0VQfRBrUKSN8ZdbE+8bry8eXlN4v2BwglSX6Ssx1+aWVvtkvtcVSPzHMo+spA
9ByMYGtaqMbwVbnQxho6ITbgx4qL68f0PuVswxQVyrtw6PEQshhYYUestMjMIjP1+ISPcOYQAFOA
q+akWGd8KWTgaVrbBtXdWXp60QQDHILRczJXkZCuQcVrF5IAp4XLUrmlcnW4Q+TmQxgM7KCAf0Xj
w+CdI/FlbiWlpjUG7OFSGbnni9ZGLPeyIpIevfZ7UQDGduQKzsE3qEVaNcencRpoXl3rT2SK6fyz
v3JjQGrqL/ikDv/UaVUAh3BOn0FXRmRmQ+MGGA/GV31VsOlVWWsInNVj1dojzdv7XF0r3Z6Uk0dP
9n7UN00wkjPfd67bRz3h/KO6vB0WaZ0tGeLW+MBVSqgh2NUgOjCEDFcNgg6NzEQnqfYq9wq9XoFH
8Tj5KfMxZt1tcf7un/wpWRlUYXhIBaiQgW8JLODUpqmBYJ429cT/TEEbxG8xXT4Gi8j924wLy+sh
rdeU7oUnSj2+jw0J23OVA6t/QBx+olFwFIl3/divsDKjtmBH6Bc9+ynSQPRygKzLz20SMxlobNqF
CNZ6rFxQaKoXbb8Qk5K7wFx106ZUvUlxz++P1Dy60uSdBahUSgy8qVp03grNoGxx10iyKxt54kXz
GJD0qwyy4fID+TCUH8SQ8J+d7TF+zNJ0aMlw2H0LvtTw8txchY04yCk69HC0JubI9NRnhMIyZYfs
LgegTRDcyRkfn8exK+wPXCfpjVJP+fEUaH4inVd46iLLM/nDwCW4ZMT041+mpSuXy44MLcxey8a9
FseUA3HL3+jEK7b1PNFgmMQCyjWXoY0qKlWzE7HUEszOgkdWkfkASYabyvANTf0UxK4AHK8MYiSm
RnqHCUV9uO7MCWcGvMd99CiT7PfYDXnYwqy+WjPUFOgihqvPC2tovPdacMIzcTNq4Q1L5lCipUo0
VzqMVtNh4ZXHwdjIgvLnGECDZVII+P/rpFcRmKs21WM5rHW7heA7754WKZV+AAcmrXH3QPYzS8ia
JF6EciXhEPQzrmGdnXfR7QoynOTchDwVPLsNQkTPXlxLDz4k5wvS+m0MNH+tzS6U2L6PP3njVoYv
4qJFK3ChxQWRIt5MWRd1cuDLMNIb5KAZRBx+g5cx1ETyUYyaMc+p9df5So4O6zG+dqchXRl5R1pT
jnIY4Lx9oWurtMxe/arWEPDI4CloU5eOAZeRKy0mff4l71Hv1joR8PSR9Y2LH7JBnxagwZ5DR2Wl
+Oe5hXk/qFxLa+POIXSwGqE+DfQKHcgmGyoaMcOSEa05X/GB1/wLahMPohd+NHu9mkZ3WYp1rXwi
R4nRvAlcZyY5Hu9sRJ0/IC4N9xrgY4i2AgRHZ+i+olrzSqS1nF+7W1toKmsN3NWoY7HDnRC3RGMt
PVHcbDwszSHySIhfpPy3X8GNGx8oBivknJJkytWtJREUdv5U+il2jdyWWKHsL8nwVJFPWNsIYxur
rppjtHX5DeS2RbWgDlOH8sxWhy+KcZ6vGej/hsEVS7BsmzIaAsz9XQQNL47dOFfhDurZbksCusJf
vitgs64MgaxQmzpMxYfKR+aHdZGl3Inno0nop1Cna5Cgzf+aldQtsL70ctx98+vdH/Z2ckLqlyxV
y+GNpwseJ5wZAjMApQLIIJmcNEO4ICggBSPDeCRO7pCbVUrj7ROqSgkoBRE/tzlAJ3KLxBiKEmxU
rJNjXDg0CQ36uQ4X/8gWtCPTaZOFDYBChgTG8B//btwfY+nptmBr+q+SvrXd5kAk8jAuM8QM+RBa
rC9AKMdqxZQ9dCSUYzNaGPBEBvek24drhT3yVd3249SFUNhOMjz8JuSmVJGo4B8XVPV9ca7Kg9Xu
gVOAQ4DxUcDtX7nnaZe5lrYjVYSDrxfkZKeqPcvSbfQUXn6qwr499w5fTton8MczdK1g1GyZ8S5J
9F+4eoZv04hAzvDwV6j7js5rAAHzSh+hkyNJFK3VyOlJ/OIpZKjtP79nxPEi36khspQPiQbZDsXr
45KyJ4r81VDvZlcr1BiFaItVRo9nz507PMpx+PQQqJJqFHQhRCDC97OwbuX4BTmT37fKnlYXEBvF
SlVGurWdwaFe3EyIPusIBsWczD/VhairAr60556mNf1SSi42C7pqfdwUEKlS+gH1hpU/weYat+N3
FzeBWTfhfveXAmZzi4ehNDmXiRGWwCWlL/aHji7HUprZ3aVSQHIZLDgCUf/+3FcW3M0pcQERkA71
/DxhWaf/MZQ94B173Q3+l9AStyTUZgUSzFX3W0Y7z0N/alZ9SRdWuwMp9GoHX74EGZqGlxeHfwy8
Kt1qOx33b8x5cMJnMif3Ja8pqfjp82vt4BB6ZPuMxygOta0kf0tCU/A5T99uPmryf4Sjfvqb9uEm
JrMvSBDTV/wmU8+QEMQ3YUrtyBXweiJhq5jWPIYQ/oTycUNUw5pN39ud/SqsIYOFGrSQULkqG+2X
7SE6mF8IbByLTnoWA0H7MK76bhJkHanxrPw2iiFrFzSylRjXSf8DA+gkJ1ZGH15LC+tatibK2i/x
abXY/ne2Yl+Oskx6iVIwhrR7flkiUyh3/S847VP9jHA9mnJ13KerAoG0IqmGAQe5CL9x452Dcsuw
sy4KkQwivbKl/r+24bTSrUg5wVjSIOXgu8aIOEt/l/jOc8FfxxcFLuHZ1vjRrScYUfX3Uh64Ok9a
dF2W60CuVC+Atkhx263f/MaWYEcapwzEkTX2wGQajHSZIrZOPuVbVW8g8lovMrEaTELkShF038J9
rtQ2oj7WKxIJXCug4kQR3awy1S0mvfnnCftWo39dTHRvpBR7pwqkwNX4uiF+zbXw5teUzzEv3Gzc
zH/G88/uFuWQw3VwqiiPrTHidxR6m2kHhdDVOSgF7i5ogRynT2gNEA3eBHIh6QLPBVu/4BO0YnzA
O1zJRMurq8rFyL0Uk7jt/6d3qD5UXCI5ymmbge6G7P+3CQNMtolem4PsUSE4fkCf16fLFII49k1x
iazLbJy0CYN4LZtS4I+/h4hiXWXyaM778BtIafznJi9zXsjTYzDXNHzI12b/czCYXB/9SmHmz8ZS
dFT617vTwb0R/EAr6dhnnVMoWz1BfGTBjc2ENfc7aIHmUfxezWz+7Y5FSQzg51VsqCv7KbL6VuxK
2XNf4eXIbHvH//rz2fH5mY6do5y9J5Ylp+GLrbeVEU4W0ERc7ljxff32t7ZIWfhMb2qJQ6Eu5p+V
neo8bNjDe0fbtj7BVUaOyRPd5nfUBWYLC40K9ghtbauPKNRuKk75JeXwVxh/bxjI9IXP264gWODL
cyf/NO/y+MSt8S6qr8OdnxhgtXBvT+GzoFq6IJOtL6yTZGVL/1ibNc7B+JWVwBAMoUMou6w/jfGq
ZPqlRHH7eHskUDsil88wQJO/hKq9X7pBQ79v3eR2F5Mwwu9LO7/x8XBNl4aPNf8K/gL6E7YBo9YB
GOBwUtmPkjYitoA7uAdBlWJZofrvaCUXvHXMwdqIKQ7U5X9c03/IUWlCWlY6qdvtApgHMxS1fJ70
gXD5s9nOzk3UwwoxzYeUQCm1s0AnC68T9675CSLTZE+inSDHz9jfNOEW8dvvSsVe+tt3V54dnXsp
tb21/kw9wl/nOoMFJo4yziatOOiCb94sD7BClA1xkX/aN3xCCAe5l7BH0xQUp4ujQ8mkADetcV0M
TBEJH9kMyaaAiOmiYr6OvaHKvmjMLMWCYkbgitqQA8pE3hV1WRH9Nvz4kYIgaD9CjQxqizt/O0TH
E55y/9cywT686q+Zz4NkFcTSugSwrg/8gUWAPuDQrT3CrjZuu3Zf1vuWLzZhi+/U0+7evLUXV7ek
IJzWRAQWAZFtvPCRup6wGG8jsI5szPxft/zWnMXXdDXfUoL9GjDgZtO3g/jLShIReyg2AiNQnX52
jA9snDAvBU6m8AC+jvlTxTEp0NcJYlntemxEitjbLWTIJ1rIYZvRIuAcGomn8Hv1+hTrK8YXOhZs
XxJYIha8fPxhY5lc2uIROAvxid1aUNlIh8VXpDONflva08aYEwwgQR+qrw9eBc1aLBw++F0j4hy3
kN2jU1Lt94n4GPdymFYNsVWYCbhU0rz9OSFO02+Zag3VppUBx/mqnIY3VU7JOFWL6xDDceMFZG82
UWoWAW7eHMzvdGGkfoG8E+NMaPRqjAv3SherqpBNgJAjO/BCShdTgfSz0qFKUgcVp19t6BBN0O92
dycR16FGRthU8tGZizW7/kNvvT8oh3IJHLtZNJ3Y+mHWq+ZkL5SoEcJYut3aew1UmAw0Zf8vYdaS
caIhEw2idNTJvP1k90xRcVfYwQesIFjU3EmRoOzccgERiD6ndIYpJuAqip0ydhwlyN2bI6lPQ46W
bOV+tP/KUnvsnSEScMqZwnfXBB1kJFrP8XMzmhTEtAupclpXW1orxmJ5qSHFKU7DGFhrIP53fSgU
D5EE/iUnpp9a1ey0QpNsjOyzHe/FATWJtos0NtHPZMiTIpTB+Y1PG1jdghx0ZZy9J1Rhwm2i1QqP
lRhQbD8gr23AjoYjkXMWDDPinxnwEMVPYKOCCr65Vxh7rTTCaE8taoS8MbYHwadMupu4PpTQ+ALb
x2iqfzAISzfafayIISc4J0ucxnyGpRNhtqICPtkqQ+v4Y12d5jO+EFXDWhBfOf4rEfW5ZGyay7to
Xlmqf80sOErHPUuDDdwi/dUrTNhmUMEnfOjfRxOAR5gi21fInSHzgo4OGNLHTcUVd8YCPZAjXfXf
xB4sOblz+yjZvMOSTgm1GkdZGEN4xJzKRvSSo/bNuxGDiWt/hUkgDenQnm7Bw0yMnnf7Dzo9uUaa
Vz+JKAavADwdCd4Gr8zHA7eNaHB1afNG+aR7q6a9pQ1HqNJJWqHE0jxjMcRvVKKO+Vi5P/a5HLly
YvF9m2MQXA+58cOXsTOy37gar1KReP1WWQYu3C/0gr2HUSsQdQ7MplUEI/zJGrqhKvY9L1tpHiNG
Z9Y9HecFpecukf18FK2fWWTBr3NcLdSxXwV9Jf63G7jtSL4DE6ReIztoX7QgsRlYbIuJdD13gUGM
Z8rLfnIhYZSaaTrrFsBYO7CGpde7xVgGBEPEm31Uv65+l0MDHcDf7cc/p6iYrhFNgop3yme+SlEh
TnQ1VmLm/OxHjckOPYmCDZsGJbNXTmZ8qzj2eEmT0CtrOV+yuR1zFMLVp4VN2pbf3BFKr166zMDL
mbvP2ITcR0wed+UelGYs+bSvV0Hi2u9XIAZGN2S54DiryOsoltkyFQAOPQkq80Fp/ZY1oMCxaMXJ
3XlkEjmgwBvxZ/gr+Ob+j4sE16gvmos7UPf0IjdppMWNf4pb/GGDyuss6OgyLjSbh27DSLwOJ64f
+F/FGwRQdfeEd3XGGAPckaOMo6GXmLbHXoZ0RHQonJP1GYpxM244MTFNliFGB7IzI4+ijNaIS2d8
r3ELhi5wA0Nb4pVt18MHxAlzzmfGgwXPEwWMvPc+XGgdHk8l5Z+v6v8h/43oe9UklRzngRUdKDll
VJITc5+ZTAU3Rc8WAyTMIXZfReuE5ixF5Ol23BlhISabImlSxxghSsI+rXSyNvddNXVywcyAlJ4x
YVmk1lZ8UXz57xxkdvxHrnxoh2OEmGQgfCcwaz4n6N1IQbhpZYY6Qj97UC+jTi/G6Iw+ylGiaIJi
iVIAJiMb4XTwYMHwqkElRpZSWmPpndpbUW1eiC04q3OBKUNZz0FLS1Wi+fsfAvKW7XpqQyfQeW+x
VKcJcgJJXIEtpvgngg2q0MeaFVWCfAH7y8lBCkZi+nN8oSJoy4i+cImSz9F8H2Jxo4wrEO16smX3
beX7r+ACMj2QQjqAELojD8O7ol/qlb6D37S91ucm5eJJwQmMRCx2X9RZVzxSelr0GngAQJI953eT
YXEXauwoMl3N57ZYn22cGAdwHQ93G8AaKL/NeFmlf0CztYvwsK+7iR3kjLFUSuarSuhkhgWVXuJ9
RIgl5ccgT7WeOKgWitrdApGehMEc+ooBB//fFiGuwZ3+q5MwjqL0kBLgSTA9Pcy7UuOn0UFMI4Wk
318I/SnXTcJ0Ohkl0wiANy50ejdIvmvGK3LrAAWgoMZHt3lh9n5aJTnSTGlvTqyNIO7U1b9yiaEt
jKCKQvw14DnVEkcQGRtFw0AU2/AknZUIdwa/oredqSLSTqiGjgM7EKMclPJhrHGaIW0O8fgHh4/u
6oKf5+WLJPxUQdUO1raRTLAq/8WPR/7+OpWQ3jw/6Ce3azkX9JoS9TSoRAS67g6yiPv9sxFMrVUr
64uPn3Rvy5yBr53cx6ZkgT36mllbU72r6H7BiBOVhpAx0c3/6BvmCIS4eR++W5AsZHTDgsKWHjiA
P28KF3aK5+0uvyEEIwMsHeMYeUk/imekdQFqx6cMbNs5/9We+PhUVBhrdRZSgyDIkz4J87/IyM2U
tXCuptbGVrjFwFDsH1smuUylJKHRy6QGmB3Yy8snCh2V6amqntSbWeDBaH4uMI67Xoa+hKyOTY3U
vqcq8OD0JeDar9KimzLg7cW6fB5W4T2+I2qCJOALPR4ogB+q5S2gsIncXc6JRLjiUlKKmNqk6QsU
jNd+kcCiK9cJuBJTvb5ZMDclJPUSR5dVX70NyQV8wtTqGXhIwx6dQGA8ny4TP2DxNwh7KFDuehOf
LX6atI0JeeE0TaExpVF5MhLxcCjwKv4mRlUFjNCYmLzHszGQDdvpYcMV3gC37LgUTcAvPoudoLLT
pRSaAYJjemVG+gCYjQQ6Q44/upLNxdSsX+AZuxBGy9m06Y8N/Zfo1SVrIhXQc0ak1N2Kc2j6dZF6
KEjlJcBK5ATAuKc8+sWQETU5o+wfdHIbs8VDiksda1CLoldlm/qR+8RUJPESb9noMBziZZXehPBN
M8RgUrP+aPRCab2MTrjJGb7t79caPVo4fqeTaymGxl9W+8kppPWYwxQRUCdkGPtOnCW12IIxVFQb
X+U4iNyDi+Fy9uuyzjSqPrMrE1Q+77MJ4gb/nlXi332bPfQ9yiOdFtPqkCS3DSvjUpEnYjYl/1zr
7Jf4Vy0ZpzZr2a/ctqcHXqAt9sg3MckS/0+1+96os6lJ3wuMxmZUsS5Rfn9D2QdMZpmAmWlaNsOg
r0h2Js08FhvKlKQO6rPxSUxVf8NYkaiz2QVRPu4gtwOA3xtryhBvsgEANUYzI7EhmAOk/dx+1zqo
lex3NEli/t0TQDT0P7d4w3llMHYFHT6BtqwsFE2LYQTI/HoiJCR4lHJm88ujes2jr4vunkRaEmEp
Q9JapB94lfAJol1si8HiP7akbNevpcJLOnc7eSvEJff8WoU/H4Y4xSOMf6Z62qUWPZ/Mv50klkTt
qihRtKQSlMWM1JlfKxKEu4c5gc1TZK0hrot+2cYTwCEmN2yDT2lDkTwZ5jNmIb4l0GsgEC8s6eAL
buuvsxpvwbaZIspClhdHpP420kBTRmx4Sd9NZzJAD3uzESPZGUMIHH3nykxDmJ3wrg+rABv76Z5z
s76UAKEUKMI/H2GD3T4YaOrzDT8lwQNxIkq6YW0hEryshbuf9iUgdlRbzmEncTazJWXvycW2oRd4
9jHDN3S+npVABPZlgW2Coo5+p6AJt3clwa85X1fLGmIfEb39rYvgT27l+u5KymYuIzTRqlFrxdpz
J61ZHb0KRaG4D5RXOJi0F9yCKnfU7kBMfQNzuKhBNn82nn7N3fml1fwBZD15BqqqSLc8ZJUJ7c9K
vlNJUpyyC5Fmpzekk9MPa7H6Pn65e25/LvLJQwt4T+9iw+YITZcDlFibRGSSKyVJftcz+MXAWafP
bBRVmNlHOtlnYL9mThHalj4ywZn3sRGSbjdceVl9navHbcYzyxzlpMnzESuJkc0N7cO+XUUVx+/x
6zFxoJbJMpS0OfSF/OnD4m2Qqh05JqUrwMSJJ0R7HrIzYep/+nfDnzpR1X7o8ZvBo/v8LwkFiDz/
0Nw7/7kogQBbMgkxhQe5hV3DB8KyRJ5+IfF4C2TFVDgP21WGFkr5pNnuqjnA/+FvSeWmPAnvpX0f
p/TnN99tbyzeHKJgIlhsNoxxTrWCp8+2QKYvXcRhflwbRJhLWB4PFHKbtgebQJKJnMNa07a7R83F
V6A9hERhXfbNpHjiD3o+uu58Y3souvLzDdgeO01VL3p0ShXmXldtE5Bt2eAfQFje/uHXxh0I8aQ/
9tcJTwXHS1fW4WGUp1R9LKeD/puBiX9PjslhDXUNT9SvKcORW3I0SIlBrIaTIYGfnFIATPqIBQ5Z
INWms5PmKoFFNbwHWtUVQQ/0zNFPBD0IULk78QeM+OQD5QuzyYNwGKTq6NLMm4cNHVBywtOClv/L
0hLLIzgLsZPlIaElfEbt0qLD13JqiwG6arCwlG7tszDUxI5qL2rpx4o0IXciZ35wgGHKAe4HBdfA
w0e6bPZJ8KB/Fn24jNzkUoSevHBcTCtMzT1JfxpHSFLRO47/kVZYNd9XCqDrcZqSD7X8Ze3x15xs
/BFDSQ9tGDAiAaaPIkH5ydWAhWFfNG5+Vl/BdqqEqdPfsJ3SI2EapjBVcxiWFFZhbumz7rySJZ0/
7v6VAkluo/WY/Nooh8cJoE0F8+OneFDszjF7D3QyqFy2x4W+a4MTZqnDKMuWuplfp/HWAyE6Ysma
D4FKlC/LZhVW5M8q91A6yKRBdr5eudY8F+/giZk7xPY27czS8kZM/nR1C7L6Cct4aA6dHshi12+I
T1x8JkIgq+r6A+GzDet1XevJihhJiF0JIIBb9CzoFvey7SJslWy8E6IcIiP4czoHhR8q/D5Qh1EC
kDgO3c9OrjRP0hWSW/J01Uyo1VfzB69aM0l4yHe6XmIuw27R4TPy2aDyW1AFy9VXjNHfGzApXthk
MLJXZxxduL9BZfYDJVLsQ2XciXRL/1nnz8cot3wY86Br0nZ/hWszW3ndQaPmNDWmqDCzMNSuEwzY
XAw9JWS5/xlxhioA4HCqAckWfTIHQxziZBTqnt/Aa8l5d0PLPWL6l3mspXmqdtdRCfG5WaHRY0mV
LogmJwfwvLL5C1pVEfocwKUuavHqR09pEPd5uJUjogibO5ViIHdHiVVaPqBZvnaZCYJczwG82G9M
CLmAYqizbvrYKkLZ+g1d4WVldIYs+ThsUMxJa89re2nbDn3e9B5C749zxaecNxZrQnMAZADwJQp7
hgE3rfgP6hfQmeeqcJBEB0Ckw2ODVJvNWbE0iFxEuADwseOUChISLyAj0lHW7sjSU71HUHzsDtI+
9PvGZjmc9DkBKdRijvtNpFHSnN5tHE7r1u2WQRwS9w3e6xSUHXKHnUoVmWg+TzXHuAusTlo96BA6
I34imRUY9zIYGJ5gF0RPdxjOpkQBwOJnQLPBC05MGE/jHR4Hdm9Knie7IB1GWuJKtIpjSiosHMzM
lWB13X4ro56fwtEPFJpQoIRM9zZ+s4MpwIfKbebpI1kGmOV4pYarzW3a/0MKgpiGwV5X465kqe6c
r1IZuXqHHFVs0BheVX056aptqJcpp/F7GV7g/3Q/MvkE0kWBEwSXDpnv9ESQf5P65pTlyz5rfw2G
Z94pwhuNw9bSgfgnR+G2jJFDbZUb5bTOtw8N2WZBmnW2nkSjcPBNOV3dv75i9cMZfzFsGICaclew
Ga8l3Alm4sqU4l2O4NSkCtlAhUFZUbg7Pehs2VFBGK9DLj06zQmX+RRKly/OWayFgzt09M2Swy23
7SbZOPB0P6ldZIkAZA6W2rFiYrcHgHoElhHO/Gw2GzzTPh3X4+9lXc2dYvRHZFoWiahafSV9aFe9
k5cBzttDJ1PDgNJDKhidkvat/b5RniEFfUHWUZKDZVv8y+qCyvxzg8irYsITd+2CPBLtkxJ8Lxo3
UXszGZYXL7S/SUIFyqMFqxni9Xqe+tcBWM7XJD3FZtDV/liFZKpFSLT2GHorK/5Edz+G4qTmpkD1
+pH62Tm3pXOAfMq4TW7YlOKW450CcL/4l+ZwdoiiftLm9SO4H9zJLq6sOIOkMfcJ70uezIvfzoP0
U3CTChB6xwwpqPJJBW7u54HA+Ccje2QKWkbdfBWT8ugUxEfK3VbWqq8V14WTtnRIqs7OySKEWUiL
2R77j8RTsygC9pl2zNCp+fPI2fBIeZHv3x82aEJg1buovkaPVQy84voqy0X7xLPRW6V+Iw3l+T5M
vRf8MR7pzqZAIGxhxRf9ESmU1o1H1yFLJNCmpdcBCI1iCUMoiNOT6rIe/fQ6DykAFt9VjSWmDm/K
6RAsVPHcC0p0GSeUhejneSv604TbT+WCNS/ddgtxeT8MtwRwUx1weqTqz3cTPnF4jo6lHjjwGihX
MnQHNrpUgGuZelaKDCDpgFCcUYPM3Xae55tkZUngOT+8U8snQm9MN6FMAFNu/1YgF/J7mLSI00GY
1jKZjwACYexQvKU52hb/atsYs1mGRqR+nLQJ145NOKoYxcp1NmGo1OBQ0k/hXCHAK+FmN7TNurdg
e2anoYohvReP1oQEMA+Dt9lgAUX9gXzcU3aFH4g6vw5OnN1c9zdUyVKCuaCUNBrPdgxV4QObllY3
3WdyTsaXr3NB/azet/I1uCm8NGsckKYJhI/dxF0x2BE9RppJmZIZHZzvdVxhGDYcRa2bzlJSg3ah
xPbAvkRzKuX/q8dtutmgNDv1IYqjtTfXIx6wjof0fLDnFhdLhHPQT5zv1yAi116DWmL7lAh6tcwL
4+tgzurAu2H2GiSXYr1hSKLsnhemTXc+dAW4h5I4qLJNl9ZNGsgbLoSMLvSizcjzQ0vhV2UA9/Sk
b++Vck4N6S7GeZGmE/AQxuB8jjmxfq5HAysPlFDh1PRbfsIrPwLDI1MMUem6Md4RWJXrJnYSYzNW
blrpJN54fDLcZl9aV6u3mhFkjnZuIBsh9ODqZiSJ30iuchf0houRNOEKOKfTgNdBsa6kLbD8yyHA
uv27QP0HivF+oE+7l4CnIImCXT/5zeMLuwzsi30VpNygUwnwuDhbdl9P1H8ewed3GxCKoBeAgh77
6BVED49C5mgZT5+Qf9cmkHnlBnc5aAHDkzcUrml6oz2Z+3uAAPXXrC+iHe5Q5BbdEHsoa8eh4ViJ
AJJnh0rKDc8QfPVazdiwGoFbOQt13jgQW8JpaLu6HrseWSh1L9IKeXlEYteEtQrqoZfqB2eMMsG2
XIXAxtSJ2caFy8lqZ/d2mUbSX2wQARXjdukPztPHxtLLa+ywsv4zQmxKetEKz9BLGWcJJDOTG3cS
vfrrs6twbb98/S3CdgpRXK+YFAEXHAtu63WFP0GGlV/dzThCxX59LIWyDGWIfiMxVQxS5hHG41hJ
b5hyTNSwGElCHSU9rmnexwfyxLrradjmMapD7Lr+Fkvf286sdj1Bzl3dAZRwuRSGWRW8E58kTMr+
pM3uL5ilBUatI8sK10knjNUWuonoX9G5+D4UpTSeYvj2PGjrDVhrnKxVtgjz1kj7MVilJKDrC2AX
07hr1BifRgwg1kviW/f7mUb63xnuxhekjO3gE4Rl6lNT4icsnlDV6zKk4/pyf0aD+bF0aP+ZAEzw
wg19IoCJsFthAdjt+JsFal31kVvXI83abnbG3tEFGPx1VltEW5kPXmZU2khTAVsodXAGNH9k7jhw
x0u3IiinyS6UoADU4VJlrubfk/LnpTeI++q4P83VSGu138q6DavVXHT7xIOJL2oriknUdRFNCP2D
0fROGB2KLgaJCU5qc2C6PXoeMZQVeqXPKMgwS+i09jfBUdA1fvD/MGRKwYqI+jQjW9K8lXD9uMkl
ijsvhOhFEK44A5b/0qUPnz9+vyQjvzpUv6Fkl0DgqngSy2hl48ntWZrxi3cVvOOYkS+FlgC9+YvZ
YpH+OxBSMBQ7+q6TUdEnXp5RNd3Sff+y7YunEHhHgkgJ9orXHHWHYrCI1PYMUTMPgSbKsy6XBLfR
GH70D2X1RjECZOE9X34+6rfvSwUuy+UkOJ7fmTnlIJdTynVW7if8jJc/66sZtIF0sfUErVNlkdh6
PKz5nQ6jr77E+I+K7QIutRqjNrvsobHiRulBq87T+Y4E4L+y9RKlHkkU1caV/rg98CkZtMjknDGJ
hbDKZGRVVjuEV9orqV3q+UggmnpdVUBlaJt2O7Ee9VNo+pA6P/3p8JRyrxVsbFmEDzVPTkEFXM/V
LHuYVi6rc42LJkyv+s/pK5AsI6yhrqfVKf0YYkbUWzxj8eCPg8h60HfWPuz2GlKyX6bg4ZeJpyus
/KyrCv/qC8F6U1onosazJhmAdJy/VKwF9JkFVWBuVoCgtoL392Elep36ucZjl0LbqyOIrG04BK+U
P2aH/GXk7U7nUtNSl0x9QPtAaIWO30cSTG1281H1tA0tW8LyR1JFCqrXqx5u9YAW5i0nZs+RHeZl
TNwslWUo4ZHgWyg+aXRjMIUSb8/ZRhQVv7kT3zNzNKdGfSlJQBNDQYKAEsouBrh0c/kkDpo5qW5c
puQWSQv4YS8rlSWqlWVKl0DgSy/yCASEcY1vNFGIYMl0Ra72S1LyieRLygrvs8oG2ZIJqL3xP3m8
Iwc93BzZvEshyIQHs3iIzJKHqaqsvpttXQa6hzVNcXh5+uU52XftfgeoTiLEvjzmtKA1JvkebUKO
v85oI9nwLGmx+Fx8L69q3UdFw7472tYd4EZWe0U8MRunA3z1xO8fnvwhk5WB9ZyqBvr3DGsqJ2A4
wHYcqfYidstTdKJu51aWLD6Yj/+bhesTeZTbPKCF2woRh+aB6+6gVtVFt9nq4r7rOOuInYjpkFE/
H/u+L9KuTnsjFqJ2NFeWr9Frik1jw9tf8Xqpu0s4XizYwkCUpw86cY5wCNBV8HpvqB64Ake49M5s
9A5dzHhm1AKVjefQYkIJGCSJIlXV3tbkmIEl7Gv3I7Sppcy8M4OwpiYC15n2PtfqVfuMrL/+476c
DRBL5JOWSRHvbU9kfG9rnH1Det/Pc3L8kHlOCUrZdfgIOrZGG0/TnuZ3meOzOwQab9o7Iwgcc4aa
p8cUfppZycfL+DjjCUzoiAjyIfQSncCiSqNVIzZs1DbQYup5JuECtxJoQd+Yd6DFYMuZeuyobTd0
sAGMEpjo3GNF/auc9N5ofSjafisIopStGMxu9Am0IPP/s8E67578aXh6WhoL816sbiU8GdgDpobE
/19bS6VsVguE0XEvfHCWam5jIAreU1Ps9etu1Lf+wfwJzyjoucZWpOzdZWpABax5/nJN667oiCLd
O7aYZemhPQxA9yuOdawlNo6QP70OC5josG988l7oDkkx/lUVCAvGeCEupOh5zBybwsn8ctp22IxR
TCkk3lDboK4/knmDy4dsIjHN6nkq8TAHVzvDIGJfs5YJoIEjmZSxO/U7STSBk/uIjbZNORmDY/RN
N0tfTD3JOAxbqe8seStmRdxd6xWAi6pTwZZjwMGSELcTogtMZ3TfGJmur4Lsxl6jW3FXMstHr9o9
al4VTieXw0DVtYjGwM8l/hN2oMHoPpcB6IFNtJdY4fpYLDViO8ezRX1Gi5tY8TQq+COajw4oM+R2
a0fZtk+JhywTdkTtyREdJVNKdapFWZbuZIF1unvJc0Zo0v05yT/Wb7sBFo5kzTS6FSvU1sMIjlPU
TTLZGnW3nXynuxcBTFb6F13PCx3YKkizsVdN8jG4LJqz2gOOs5B6T0/yKVyTV8o7dBW5v29hpyI/
tKl9qseH/vD1XN7CCkbzdmjvXwzDwVBervq8kxrpGAQm2CCt4JRAsm+uMNn6oZAF2XXoNLMPrx5N
9A7eXi/7+I5VAgbamYnyogg8UQic51/5UdVYkxVQ8FLvE04p7CoBsXm7km9S90BChz34eMX5TQVi
DoGkCnSYjqc4Q8z82YqhmoWYvvHARH1UQhThDNl11J4yHCToO3mDi1d9uiT+vy7ShlgxYl5vIbKt
Ee3Igg2K+IIUuvsT5lNu/VS8KlgxSoAfMimUd58vPbgr00c+GMOmN6GFKZPhWk6C/w4Mts4/u8wX
wHWkxnTFu5HLybDZYdIo5pcB2ph3LxfhI7FQY5gIBIOWPiJ2HskWbQRmAcEhLFLkghb9ffOKhoJv
EFcpKS9wJFuakLaAnTJi8J0O9mxbDmzemtnugMCf8bWS/H8pfhyrpE5OR4FHd6wmw/yDOa0ym/YT
1i/a35Q+jmSEC9flVahJDzw8nlz1f7bPTt6zsxg+bQHF4Ev9Vip9bU+tpJG2LGSgejzTuh07N3Og
pG5fkpRH/cjUqNrCrukelFBy0OKGKuRiSAxMzAE3k9lS9ue5Gu4VpJ1mJeYLSKveBb2+cpDZGqEo
5Le2SVz1Y35M4La8L15Or2nPlUOmeXJUzGNWF6cY1jLZnnVJEVF63gTfI/n014CM5MQGoZ2BEgic
wMaDxQxfHt+suY0dclYcY5aQWAcRjVOfcidrsLvPz7IP+FPh87GVKvuBkvvJVbg2CT4Vsbr5PYSf
+2UGP7f/3wxDd0yUGPHD3VfCVvT8/6OP8A8eDMeND/uMF5jyigCgGI2VS9KgpbzFk4DHXpaMHFxa
Ude3DsmchligDyG3crALFuLzzNajuoz7iU1ldcdDm7P/N7t7p+/YgG4Vh0fwFC8H22GLPVZjZ3FU
IYaBDxNOzuAcG9FRpFtGwLhLMjgJ3NblGqF4RWCoQBXdsKJsOIXV/aYJJKoUT9IAhNeT9Mc72hz8
Xgbq/js5XuB1I1yeilwwg/mgMXKXdABuUX8rF4iFkVqhVwo5comnzfs1nMYaDvZjHNxwZSergSgc
WdjjVBmgE0ulDg3zXIuvvFvrkX53slxgZ3E/TtdpVT+2g1Ib5wbKBSUPXw9V+rgSdaKH64WqE51H
hILOpNcLsAd+3x+DgGbhfaPVBAKevBiomAZyoAeZvcl2B5Z+M2Tj/J++4BNhAt7PX7y3/8Y8OshG
xmuqJn0UsCh33j/c1lUgIykykFMddZyrYKxsNABA26ecD2V9za7Y5drd9dwB4b+o1cfRM5wIQ9hb
Go1TWTKTsJ10Kjto4fhn4UdQAhCJEnmkF0xgesFfTMqNdDPbXBDVSfO+l+WZMgbDDiYpEJB6G/8A
ecbFweK8AvA/sv3aZ9GXaZy/azd9dGS5gvTgw2osjIVkfY8I/zhzMhM0LlhMLrhBx7WTDb9LQ90n
bbZGATL1bU3Uf0+aLZc+MYYqPujzigxk+v3kyoaiCD7brrL7y1bmfrLmB32mO8OjoZBZETnzj1Av
fEE8HGtg8J+1Wjs2ZWNOOVXXdXXvN18TEEOdYaX+vqpSs9A8uyrfY9jevev2ZejwZoki2uq4gDbI
PEaC+zcZRTJgYHqPJukws+zutTFOsAcuzYc+mLf7M5KkJOAky4Mo8d2jFiW880x97OPiNcFanCuy
X83rL8c2LJDtLdIEnvdev6wu7KhQql/QYwWvDrNgLllKy7/Bkm/92TPvW4J0fY4wlOg1c3CXOOvn
3Hq9h0m2B1PKDzW78lD9H2PnqvYrIKnKzLQ/SI7pnMKGhYME7Ikl5T+uChKDYOqGGoWmObHucM7O
UCmYcyI4A5dYMLBYTAX2HddYM6fxHamHCzZOvwAPkfqicu0jimJZCYrzxJKe2ZKYNxKPK0eQAQa0
HXZpq+yg5YxBVz+jL9pk3J52I7rTQ5shKlPo8NLX6+m8iFNfnt2aTgautA4+oL91O3zPWJ5zRFW+
Hn5PujbQai91P8PXhd2Fw/jErV2MnnKI9mh3EkpYThrexhTJF3nWNTS4lI+hDUlCLBAe9d8mH4aU
yDJqDHWylz34XQCo6RVnMPM+FWN9eGFE9edy3LOFIbpUZg6rIZ3K5E071iCUTJZg13/fht37pmmI
ukpVPr8H2JMgbww79cuivg4qXpPloMoGaWezf96x85717FtzfwPWj2oV+lNEzO80WilCw8oIJmLC
6hMCDS0IFZiI/19Ogu6mYGiHthINsvui8RsrcSncxTh7KvI6CG+9QtN3C6gOMEOjM9w0Srs+wYc3
GqMPsefurgGbqsgDFV764Uig8+CkAXMEApmgr0O4tAp3Lz1oCZrvYzn9hW8AEXZvd09mbW2BtL//
Izf2KEFcMoq+fMUDjohZJk7/Ka9oEib1rWfm7yMt0b2lLlAwF6L+0PLFAu5apon9w15C0qcIhNtH
5q0gflOAarBhfzpM9oK9UBhVZkINSG4BV2EizLkZyE4B/h/i3PikpqZP/NAt3npV4nCSTApxVDOM
ZjHXh9+iMA0qqWTF/JaUhTOpT5Bs3SkeKvK589Cje9/PAlBWWo/0HAsQR3dMTB8utHaXMIKJdbRg
5O58ISGxNSKVsE3QCHADFnUaCuXrPF8sUCYMSVsUdLYYXVriSgOKi7wwQg57iveCmmulLd/0sMc/
pq/QRzHaMG0f+h2Jc18l1nrcCQBi0xnW9v92Y4OIp9/YS8MrgRf8h68Vdv0AmufIJweWXt7h/6ED
VFAhM4Snl0HqaiZNAKwCsgEWv3fQG07wW/AWBlnooycQYHACcFSSwGeW/2k6nnIfMCjfTHMUkZMe
8Aee+0QPbP5MTM/93Ewin+rU35vt5205+LNkWvrVc+WHX+M3sXDMj3ILy0lV6OArPH+HBe9++/ei
x6KII2Z7bGIx9xy2mMD1/7+rPbe5FtGSIAa74XDN8uSRlIDOi3duo+ihZ/+Jvzdm0+YbxQSqsWZo
2EvSMASb8SQfCq8W99o/6hehFhZKzeiT0SW7Vkhjsihu+V4BC7aTc1vFHNm6MuBvt01h/pfSUfjA
2xsM49ifZp3IgYmOgepkBEzaf8Y6e2iTtXLBVKf+IQC8pjKdYBb5NWBsduQOc7OO+BQ8XDKkgr/Q
frxrKlp4VZmQncDYJ5SwllZWGisGI18wQq1Gl806JEZKcuySowCgkfSoy+Ue8vqn5TPw8E/NY8AQ
TRNi0RDTc50hyg/UwuItyv49wcqbuJe/prkbsLl8V1Q5kWaCRQE5YvoghO1Gt2w772DMPX3ZCdgk
CH7wzR/SzynmvFN8uS47b4DcbEtgtgkpZjf3TVibxOaC+4cVJCzFdUVMEfcfwjCYRWC7G1NkMmoJ
+gshEXxvURyazxderJXkt3VN9pxqMG2ABD8zgafHumLNVjmbezpATt2L+N6oLt85p+ydpyo7RpsR
hL74OYBiFnTluh9QaSmnS5PzCchPnW4Sdq8HBoV/4fN4HOi7NKG6DfGpLoms9AqJnkwYBJu4L9Li
K7ABfUipZQVSX9q2SX60M5kiqcb8XwMKVR2kmKIrsqlWsEgvKs5ahRonyC8lnNDYvPcawz255hes
MxW+N5DiPFhOTX2N1eAAuKV6u0cPbqDlegrSIAOYfVFvsSVfFA4zC4HKU6aItJXz7UXL4ktYR92+
hMpBe+AWjCtCrtu7NuacWZyGsTmTatOHZTj+7tJRNhoCgocEmk+4zCm1Cwfp3Jaw8NmLNMzynVxG
Lfj42wX+w0x8AfbQL9B5zKB/ZMLa5NO8PoBFKwcAXbmUQ/GeI6igH/xVvMJ2AYIHxdK0dP6G5hLE
Wi84Ib1+9IKEoD6wqSlJKIfRPkoh77ku40dkALzksCNrymar/4qlrINjVMYxS5PSD5MCz2+J/wbv
zCcQj8kAfLNYdI7rIuucGTDbu6svKKyPxNHIZcuZmX2Qv/GvEqQzSYr9jeNzHuWWc899sHLwP7HY
mzcDbZ04MCtjEanwI2Dsr2h+Ud9K0VJ5lclhH85L90Xq1DYSb8qqbfRPc7nIFqRnQEy5qZ72Ppor
S3U2i9czffTh/PSFbmayZeVrRh7GnTJ+eHR1yKgHVN8wO7WzkUpbvq1EBlujI+lDhMD5RRGKIS1Y
sgMsKpWNWCILtI6HTxuJkEjhx6zWQRqr053vr3q8Vx6nn8e9RSp5nvkUVehsroU4MrSdDzwh1dQL
AwWQr+53ZXn8cY61qkGlzKY2NzWePG3RK1pbWyZpWILONfjWlX9y679CwGTOAJw4ed3eBdaWL0gG
eSIXEzKHyIe0oY2pgNd3VvB0qDWLyfM7Tgr1aKVHOQ9COLGeLRH603IAHnBlNY0tGRmJIv8jK2eu
Oz5siiLf0ISZHEt13NCUeBDfi+nGGSqrsDCB3Vr3wupACbhIztTOVsJLt1WSMlup041YUcsExDcB
IBPdNrmDKGQzDLhdOf5xdovQBYoz63p4PC6yGQOWRF4LzJtz3mdgWzJMZ4wIjG/p/TFujJ/E0Sul
Nv4v+8DhLzI/bfOM/h2ShmY/OZ34TXk1q+UFXwsbiSnDZYaAtKkL99ykC50Jm55vXbhdZuRPLTMe
KHKcr7Yc2ZYPSkiwXUJBNbLiAkLJN6kwEFBdLmIqL3J3HDRiOO4EWxmrJvQavbA4heaCjx0347uY
YG1mAS0/qfFll9VhR+e/4Mznw2NnDIhaY8jly3gTf9cXuL6a7tM8PlIXHFMITAfPxQ4QPWHcJctf
WfMgUN8/V4abthzP/Oo961GSFHe9dnzlrH1iunk18HV2HoQ18lpx5Vy0Hqh5if/MR8vTk/dzir/3
qetVl55zqavDnyQXn4Ute83WQ7XO7LckeiV26y6j5kJrF+TGKHN1sv798IhQvwjdHsieC1tnGoNT
ogAzgoYjUtxnQhpk/CLUBuFrAsnfKSAM4zYNoTBhdshnnrH4R6ilWrxgj13lzySlVA735EWkKl2d
TBFSMefzdCsuRgNPg6jHfO5SvkBTrlmXeVRAzthzzkYT2MwHI3lIsoMlPollZaIXuTvxRSrULpSR
p0/j7ukqeKMSZePaFgq3640LQYEVtdloduou+blFEVCnjp3P6L9dJDLeOdohhL2K8RmFrgxwRp34
aWVuMk3B90JTXkPpk0NoacDaE3qTmAs+Xc1MwTmaO4tfVwNJreJt7U16qOw+86R6xCqKfxHmeVdK
Bao9LUlpDJW2UuZ+SViZUJ2zdc+pmuENbUUrK+cAnkGfqulJoN203xgE/Ej6SKl/UNeiDlWQC9pz
47iyXFU+zGGFOc6OXe0dS98ve52Ih/y8nMxIZKjJmKiG5u4/ni3JUBQtbvJdNtDMRQdY4CS8E1dz
+rSJlv+j7Corj0KzwZVL131t5NBRsRROz828dQHxlUAVIq/DkEeeccB8V6krKwxtp3W/JOqCZ8Y1
PRNTKvz8kp6uTtsCPLuRNbD/siL7RwY8WhUguakVwrvJTmH6rKRvtrrWDZDEKYhclhxG2kpRkvy0
0rd/9FCK5b9RU8UQk0CD5ixz8ivzvz/PihKA6/bFkJDxqFEvqCwpWVNHoi3JnuXuNyvKYLETUVSu
gXiGBG2NgvNf+TWizgn+xt6R36L8v1oY+bBAsMWFrA3CYyTBxqScCs1oaqHKsJGDUiyAMIf89YHa
eZADi5ZMam3R22Gw74bncMGcJ9mgTXuWDC0DJw64FMaL4xzPjiXQn8RRQY73RA1RC+JDLBKgk41n
vXsyK6yJjMbqBsG27PC1yDSwL4qWrK8/kE3WoH1RTmDYamOVrNkq0uSL5xrNnr5p8ucfOGXq8SsX
x9vpJ8SDiPVOYOpN6sdpc9EpZdFTpTcfreLCVUdkD1Ewz4epXXzxObnXEUryXECzsS3nx2Iw+yYz
8cr1XZrg4fuVlrJjiBDReJ+r5JRfYvUWBUAUugJIZpZzLGlVteluPIN+I+L6t6IEu91oVvilbWV4
YhBWD2gqnmD9JpDXIUZK56vIEUkVRFqE3Cs4ihI1lPzuYGGnHB6lwqThuJntEOekG878hw2O/Zv/
fQIIOiaD4VhpnemyEBKM1gGILVLGMvgQktsJqVl54wP90woFkiJo2sbDheroa8rF2iiNT34Hr7/D
Mis+maU2XBU54ec8KyNYoMR5LxtJgGbpiCGKD0Z64fMvsVXLOfdRwqccCz8c5a/e2WecAs4UN/HK
NylF1UOR/MQUp7wRBxyz4qfeW9HPgl6hVJoOshXq0YCCOUXjsQ9nNf0136u5ReRkOCupyXR88LoC
+epOYu6t2DiK+SxeDnZX0DtJWwpTlwZc//CmmuYAMSYswgPGjb5UcaJIgInRRMiAsAOkFcrZcC2L
iqkMiV2fkXHQJbQMPeOe0YRYor7LYicj2wdypfddNeRhMI32674ixXj4p+CMpL2euGKEtn1oI9iH
xNQGYmmZEqPPivF6uMlTq+oOnfgZvqPakY8J8NQayvS8vBuUWgjpo3O4hzUOUeW/03j4QQkyNndF
/ortFS0w1bGpSyWbz5ZMoE3XZyXQr9EHSKZMBvSC6P089wp0EpFwX4vFULxg9cq5DE04WqGCmfUD
DtIE3O0+dQKUfCZcMRf+naDfin12kLKWP45t3babBAH4b9gPzreppvuaT2F1ESE4HuTKlBV1XmC6
uViDvvup5xb/agHrz9vYcM+Kk5ntDHp85s3swVZQMlAcyjl6TFqBdxsdwFgNKgLL0Fgx7BswVyUH
XXqm/Rd74pvnIfg1Xyn+1rTyA2g2c/7tujaD8155h/W1EFtQvSXRcJz0aT7+HmJm9dZnj4jfF09B
ZvW5TUbZn63DRvBG1+psxeXuUEdigMn0eCMAHNb91fBOsNy6XMyotd52v+Ed8rvbRuME3BZYO1Ih
2AdrYnz53NorzEH35rjxlPynBYE2oioUtcGZwDbcuLfrpLGaAJ2vOzQKq4rQOv0w6lgdgpHcu3wY
alvtF2ZjR5HGtpT7mGDZgxWrqi/j+yBHCOsKcspqXipAAgEQl0vQ4LdWbYEuOPibYBXAI2qDrLI3
ePMf2s2UQQYmvtOip2+d13ETgdZHGY02Ibd3dWOsD3FrqcNN2+jUXauLUrOsebvaHsOP4fjosto8
X1E9IeCAWE8JBvcIOTDTlJIjBUJp9YSVzA43jJ2/A5oV5k3hZglrTpQzTmZTft5gXhekGNur7jKR
/9F/3RfWdbgh48q1/KAjfs2AftnwrUYXvzBR6+zE0T0CBHHkNw7+kLp0SlfN6JMZHJLvtwXsgFJ+
w/GFsYa/XHk5clWSjjSekjSvBaB7RfcBwoIu89mhVXDXusVT4XLmfu2E5mRMvL2raQpRyX5hijje
hnUrBGDWQ+r6MrjhLM8UFtl9ECtUpAOSbfjInO8U5FKfg54Mv3EJzuc6umMgsMObD0XmyQZfBg4d
0DixxzfEoPhqKIrisJOi4pX+o6luJxRpb7NUQtNwikQgx23kNPoEi3ybCqzLA69d9mv9i4g1rKYU
YxcdSuwYxrkR+eYzizKhIeGxeaBsvumdIgVrQbbhXF5z0RxMQFuy6tHC90gXEBom0mqllFfFUfg3
o6e7CmTxES3H8vNcQ+aGYPK+PA6ViDTD9As+79gvCYrDy6c3cUTUXl4H4If6rzGZB3qkggmbroIR
kk4AsMnGgO52QjaRrSet7DS316iKjALOSObXO83kVS6fqt9d1CKCKYqcRYrrHExs9ah6cuvalxhI
v7ce1sK4UUG8hxYmBi5bdkvnEXW0lRiCiPQh+cbPETqE1fyol7qAsdjh8gIikCfxuu7KwjW9uY53
NSXwYLKnSB2WfjTtXeiSNvqbT1TpnshcAMEJBxHLJK1DORsUFIU8F3rtviGlnpf8uTNDXOK2my2Q
C7eD72tRKjwQnpEu8iqFxhLUYU5NboVlRrvzojxYs8amyrANpuEAlgFnRSB/WgbUCLlrfYJHfoRd
rpw0ikm2lVJ2MycugOITkvqnoQJPunNoT1F1fUUHR1Znm+rrujJvHIlRaWBnI0vR6SFBHMAd4qNG
sJ0MV3+ip3rELIz6CgFrc2e3oT4OFivh161UfJw5xa2yJXFqPxc8HIA61aGZxIPecxmEMrUVOsa3
lHdJRVU6izNBvUrmyj28Gu8uui7UKEIhfnXOBoRKdA2enkz/qHVWgaLn9tLcp9DOZnm+zJR1b/wZ
0OSWo6F0/fKhUJpnv+WSJtIYtgnS5WfGOMJEuHkJEz9CFehTXYnahdl0Y2qATPRpLInUOK/d2WE9
sUA+cAEKs7znGpq2OJmAwgK94pYzeJxK1b7mIthIzpIomQOBOZSRAu6VecrRCQovSDsQWudCqXAz
GEtkM036eNcBlfpoxqqFtZpMlkfQYHi4s75wHyWU36mr+IoEujZx2EAE7Qz6VOj0k2sDPn6sMmC2
C0fnfZyo+xiXYj8seN9kWlEliBi9c6EXOnsJDTzTH5aCAbBpdo+2L50V5WL+Nad7NiS6U+HFxvXD
ctX8U9DXFiWO4hFtJ0RVY60B9pt6GQAyRq9I20+fmaknE9gbFN9Ybyc6cEWQ3vZGaa2m4Jo/+D2r
aKJ4eaZZd97PgTRwiNMlSSQtCVAEpDLO5YDImMmMTWjYkh4Gos5koYQCbWLrB/ZSbbioThEoc0EE
hbqevL6sLI3lJHPQK8ii55XnLKvMbQ5tFrp33OJzVSYxYqzjNRCz59CKhd683sTZQuroptfuf+ji
9CW0RLNnySRItku4W3yU1UPI/6j98k2k2s90iZp4o9rC0dNDbc/FjcsIkhKIV/ZTUSz9BSRhlkVo
bexIMWLnV6ePyjR1LqPpozfI00O2GaDKnesVZWLDk0rsVkklpvBEESkc2mVZ1xuHZw4poae1hcyl
Tg8VaOkw3Xt46AIGCjB75I6si9LhEwXA68a95SXq4tIafuaZHGOOziQRRrvgHSI+BNtJV8U1fExu
706dDistQfBL9p4vnOeWATgcspyNfBBHTNPluUcK+6zVE3Od2hYpvhv0lP+t3sumOYUU8tL8b/1B
dMvPyqjs9Hy5Jh0ia/N+DjB/LkHMhG0pmIyOK23K2WmWxT6WzlNnok4YwEe83DicbrnigZC7HfC8
i+YhvAEAwM35AGhVvtv90/qypgxlQ5llTlvuQNI1CAKKw6wQJrsm9CfRxg9pS2SVscIkEeGA3UYe
0THgyZ6lSqPBssZ/SIx7HTRowV7pgz9O1G+/OqZKPNUQ+eeZmaYszEWSScmQxU9FLZAzUXeOIUF3
kehLAgZVPB7InZeG52GweZa7D+ylmMbMnFMCEQPZ0sNBqh+tSz6mCfuIL6PwTNTcHk1lRhKJ6zJb
bWWD/AoI9CW15VVGXECOO35FlEWdb/iUndCI52RLrTzu7x+taGHPhxHiu76UEZoZjcPAfoK8sAIF
2Pn5bZL7A3SAydwuP/Imdp5WSXCZjDzWTirMJVE+rQe9fY2LDlrAqS4SayOEFkuOVzjHWtJgfSIC
5dGiU3x8Uw2JyHtU0cBtsS6NUTrTnJNOSmXrz/vpsVlfOF6VzmbqaK2ebW04/fmVB1VE8k3xQbxH
aJFGk03SwwSeV36wQVRaCg2cQWwlhvQ7iBNYFP0SvsMOOqmk8L0ufwxGfAGfF2Qi0zkKbpBB/9qX
yxQWCVUCrsBhknPG8JIyC0Q/P1jhdgCzyy9PeXPQHT8PMlB9fAEpJ2xTr/SrSmoS++NFfmNn8rOZ
2YAFdGnV4m9chxbl4c0DtlSQQk7g7QbeQCH+4X0ABciHIBWclX8km3QlKKVZZVx71jw5Yj29yosP
Bfn0EzLA8/2dhRnLyEDjY13+gw3tFK07RllayHiBa1IyNbgAKMFGmAg0/FRGDRpyIJSN7jFmORP6
2b7BKI84dB6WLLty/v4ksBUwl7GhmAqHJsrdlam44DDwgF4SLnId9J0VsRa6L9TfILHb+bhIPwEs
MXv+lq4vhVCjb9NhF/5q7dXGCKv5PhlyNhetMT0PfuePHGalHDWFmjZ1CTAvyKkJjs5uI1JBrK/l
FwFvaKsdi5ASk1yxtKMzIGGGncSoNBORFlc4o91lCOrn+mM8jsJNWrTBv9IHm+tTYz0JEW+i4h+9
dGmNzBqLc8NVkYfWS5u5hjc6hLiq6ZqGgXy4H+4a2EN8Xl9aUZ9SdF3Sl+ek2IXi4EFxPuDo1fht
VuCIlxgBtFHBzdaF81qRol3NLQd2r1TNDyJbsgJz178XjLADB+tSZlojtEnHXrLHan8z41s9u98R
cdf5kTiwvFJuuhUROTgz6igQekAI4+nnfB1sG8a8wS1a2dARaoqVkmHAJnWOip+pyitBpdCW8gVH
fXGcHVHuZYN8Vqoml49y9q6HLrkCY/DnuIr0Az87QxbGoM4a8uIbPRy2j22xR7JOzEkYivjSyhUn
ee6pBR8/R8YsoKGSwuJaOCawkvQC/T+7sQzILPjCJo4HeTpfeip/9naZqjfoUJ7QSjj4hB8+NsX9
GXdOUY+ihByxZRhv9o+UlXNyqHXlBDiDEBSoVVsyV2azsh8Qy+knKTBVqquJEUfAGjERSm+alfYP
MuY+FIYIIQKELFb1/Ktly6BCUr9vTHEqgbJ1V+aqwBSDcsGqN9ecicVhDinzNJsPcn1gM1kMjogK
Y1Z4Q648/JxKlVmLsTasC2xzs+yHfI7TXhuOyJBxsMzch6VL+3dJ6kxiKzskflAoaNU79YOB9lkH
ND8FUnwNo7IaNbpq5jrNQ17CL9WBPtfNnIcN/i/3griQ4DFswDDtGlcyAidpswafHpbDFyuciBQr
uma39FcIQ4ZY0TvXU+QR3wrRalOM/51Vla+c9WSzzCFN5QSx+/aE3AgwkhJ0J2oun5bjZIVM3cbH
B1kaeih3tdFSAwn0q78SYlrzLJIZKtxGgVZo6e8QdEoMT+uVJ16GjlYQvbJ2QcJ/U4HSpzOOldYJ
WcmkBSjOXaUVVubcAPlwxUvKFBKRhuAbtzDDgbToRRwyC9kwGCNttve9j3n5nmwTP3H9S3FP3/F5
+3eFc7WOc1tcw1GG1wvTPCRJ2pU6p9bq2ye21vE1ujQH7f1vEXFBTs3ubqOh458/xjoq50jOhOlN
TQh/McDPMtcuHJa7f1O15l5aAM2U3pwHlxjhmuSCXPc+Bm7p5VqG1FH9n1ds25HxZFS0+e4uHj+m
RzdehW52vrwCVLSlRCMW/1Kxzq0fw9P6zazNfb9Fg8Rq/k18Ex5iS30UGtKxeQCAyJA7NsrF6hju
nhuWFA0hNbUiyrjBtcxIznpNkbzibpk7msYxrYSBDzSMTkk0h5J+hJPAbTUcVtHAMN/vQnoF03th
INdqmmeeVHXvI3fSrkAP9odhc4R1/X3cDdsEe3qa8uquVM6YUL3YC+TIsB/b4564ssolxarSfdep
G8nTLxIt7sb6+wDvxV5i8b3o9F6iW2oQ6BO3P/wS5gvNVUPXFSCTIGKhSZHXJn4JBRsHC9Z6Iu2o
rSxB70iDfU1MVuog1Yvfwr9hmHHAmL0WPXKWSaRQ2yDQFNJfecF6jP6irO8RbsdLTzLuU9yDhfPI
gB+YFrQewU84eXweRD7QUFx65fhHWBJgcHZyqRxeSMj081s2F83HEwgDUkqzV0d/X0bBYsBxKTBY
Vyh+L8hIJoxV5422XoxLNU3mRmsms2EHJY2JqodcMNkKtVtxrpXTxL6yaUBRzVs5gpffB54s/TVq
gz0Rp7lH/LE65zHbc1vZbj5bt0RAShC0l/5SinYKRFBgaKRujnsBqeU3Ud1qfnNax3DH2bwT7lEH
hlQRhrE4YegB5CmLWD0U3QisW09OwV6zArDPj0tT9ADptMei5P8sn1X6K5Mo3b8SpD+v5ynWZx7c
s4TiwM1aBA40VQZKAX+c3ZHcfrGTyEaO5VsVamfs+Mw6zn0/miW2EqDe68TkqNAzyA0e6xL3w5rf
EBZA9xG9tV9KnVBz7SRTZH/B88LLRzd5+2okrGyCnQ2wQ+JilvJrIYBmi0P78WeaLhdakpwLpQMD
kBT++RojA416vtt8uEE5WKxTAeJlWVIlsGwzmcAFoo1ohkXbVXJUJy3352bpyn1g1t0xodoV6mN6
MR1PhRCoyxw6Gw136bef6813Mi8o3CGSZX8Z55/7jIdUU2NbAiQ4JmoBQVAjw+vPQyHbhRK7xiq+
FrSaf/AT3AReTgtwRZs3kskKVshvfc/EwLBML21CO+7jsF2gzgFBuxzNqmzWOkHEFcNgFVCf6jSu
29NPV3iUPsoeMDhXsHVZRCZCJdVUf/u7D0CrLocQhRUH59i9QWIHEBBS0XhLE8Nswk/gRoR7CTUr
MXvgYKw8bsLaX1dmVrSfjOoycV/xC5OOEo+k2Lbca9ku0TXBolef5uUUKa58uO8wlfz/SUNCnBRf
D18PtaMQ9hAUNx4rh4SVSlG4AFh14o58EhOOVKlNFry38kzVAMkeC7CRc+ok56W2AIpJZEwzz5Zw
SK9k1IaWOFUWJHLbBKWTgBgzH2epE4yNqaHULQjee86VlJNkmmLpCWIYVHP1CDKmPxwXqF9mLa74
i47TKxkXy2Ydbd1gcpS1SWZCPDW6y1cB7ibijkKiJ+mEU4F68jYvXfdGHUl6cofj++rztBS3RGM2
2bRc+a5bmksRpV0sTlOZae/UaVlI5SDtLzKcI7D1SztDU4ej2are6Uydi8N2Gyb7ckwAE1nckKTS
HLOXoC6hYlMI4lHX8Yp28eVyVTjg1ycZbFokLAAk5wjf09auYdyjimycHuaP4Pd6uJeYeejNv/SC
KoHaOGIckx0API34K1VoJbWcijOitZMKWFqFmacqbiLt0QSztrDNlpyZ6YPX8U/SLDg5JkBDFFQc
D6VoDStSubrcWLQX8UNBLxBBpHganFfKNghmhZCD0/OF2PVHEMvKlT+inqeB+scrTQZ+lLHqLnXu
aGJTt5vzfyrkSBW1orIb4cNwTYNNlPlH2ftYQxF/ZiGsiM69NHVCW9GRyahTonelXxeW7NiACD36
pTOOkkv/joD1lBbhQGw52+e5AYp7h3HHNMYmaTB2PT4/KOHvA5pAvtFjHiPHtfQnStIyxkNWprRZ
ZIfkX904T3DHBsePYdFl6N5EqW4c/6WH/S9CAs5sDWCvd/Gll4VuZUTMLPmZJQyFlccs5qfEXbXT
T1Ys6nrtMoF0STz7m3L/nMXGbR7v37sycrooqzR7h+urdDP1CvsqiVIKPwwjJD2I3XhpQxZ5DO2w
zOl9NxJWXeS6C05m5XX1k30uJQrj+d4hYMxwYJiUF1zWKnKcr2JjDhxYmZtlDYqaglzhm+qvY/31
rlOR1SRZDei8w3+M2DQLLHpWJ62e0vtOpZccasZzgdHtS9Cs6GwidH51I1tnQH6MnCxKVw90I0l0
HS3ZkA+BnL9qfajU/9m5nysWGjA/HZ4JY/fCrmV9Ym6P1FlOjQq57aPcMboDrFSvwiqPslejCL57
ucRTPsfSaW80Jt8UUHAg7Gw3hgRipX9LjnNoJOFmkhKaS4nkw6c6ZyXQ80E4ll1otsZwIsI3yvTx
QBEtC9qCgDo0+/cmvMLxJ5fxAvcavuxohUWGNRXq4CHskv0uru/VPApR8n+q8NzfNvrCzbwiIYmj
LFHrGLOH9MxNhG5Ztb9a807gO6ao4B0q0LUGP8zjNdRdQ3ZlG2CUc3hujK2w7VrJgdSs6UdCG7a3
BIx41jmcJeU8zTJxvZbQ+FdAAVVfEeV0gk969skjSTbCFFofEyim85ZpefW63cxm+ywDbQPRytYW
4ii3FpHLmMUUKcuRo2S8ootC6MhBOuI/mb4kHsBDtCD2AK3lsyNdOg6SDG4wgGWHIVhsx0jKwuX9
Ze/Iy8BfVp4qP0QimT66d0gVURW8ugQPYf7bcw3y1I7CEany0ISlC+2CEIbRGw1YI3+UFyT7EwLI
vX7CdEVcroKymtJlXMDT5tGu3M6FVr3OS/yYDuTNtsxkFDNUIMOO9yEXLtKnMg+UT+Sd5pfCkLIl
vZKmL4ato8LBI3OjaEHeAvEPA44N9q2D2NWp3qWrFuzdmo0oU47d/rzAS/TuzD4ANj9KpJ7TjN10
eRgwghNnPxGr+75ZkJaCGvtLJBcmfokn0RNT2ChHk+A96GWfvvq8jmuHKroeeqeVCBrmEeS8gx0c
Th660JEQDnRYF1CoqwKxuN0ibOd9Kpsn4FiNCWBBxblnw0Q7oOfs6jWHfNLB/tohBGVn7CXbSdit
hKszDKnkFVLAq6m0/r3I777USju6iiaZWm7GgAC2Jl4qjWCuBe+GGQC7k1c0rOGw48YFF88Xj8Hu
0J6Xu3l8cDERn+F3qr6h6DABHPydYOCSihhYyYI3EyrOiM3ttxEXYUQgm9vwqXXs7Nq4qRblDVWs
4DHdM+khusm2gaD9dx9pEDGalE/RkW+DKwD7huQ2eaS2pvwgiC3Aiigcb3fzD2SC+olez03kWPHy
tdyGAQIZIC7dJax674wQgArLXQOjjkL0qF8dI0xDQebX1WWnrn4omo5SYq2GqBXkrN2LovHW2nuU
OxKG10jZ9+KhN+le2COIbkuT0bG5NJfB4mQ5wyqeGzeqfOAL14pEO6KeikmzocaXuTpnsvXy3vVx
WWeZRpyLM+IrjhSkVLR0Whm8h2Vz8Gg4U/C8yu7JyRwRftKNsVhdl6eNnk0cNuaNM0V9u8pEmTIw
/Qjjt4cPJz0S6lmt72N02Ju0Q4j+T0JqKGynTHG9oFVJ+XFvx9I41uZGDrlJkHnYDQjz8Kxz9ccR
Hog29ubYmcmZkrqeJhINmc0IFvyyXsoQI8GX5gN526limE6pfmixW3KnZNIa2Xxpyx/22vpXcu4k
95EQfO777RIPFUGS1TfnMaTe5RrZTClsMnK9CVq7XygxnQHVVcf+XqnIupAmQjy4qbaTCOlg8aaK
Y1T9ogKTFRL+7ZTId/YVKivXjA+t2K11+ueJ5XuUEdAKiHXPs/HI0AUL0VeufkVY+SETQJ+0Vlbc
0tbQHKjn5pv9Gyu1mrkneGqzIocg3XyC0ZJdiX04yG1JnXgl059w1oSWbBx3R6RUgpbKiFpiiUiz
jIU10mRaZBahk+ifEzPJ+trQwpS5mtSyauuL6vEOYA0Z+RmQwILfGfBuiVBfw8fcwbjigwKtyxwP
5c0mCeHcf96fjxVL9RGhwM/yb8lw1pn3ElF82DApUBSU4zETZhURbrL3hj+8tdY6Odyd/juGFZXx
1Ia6G09BqC17DoEInzAeGzwUSI+IcGiShlBc/kL/2cUDvgUoORwVmbPda9PMk4pqj8Y5JeFafABQ
Tw4tCfEZKXKVmAWCATFY15EStCKPkc39OGLWzF2mDdybBr7lctvSQmKG/lJOa3Ta308dzBxQHkwe
eBJxjKMMge5y83Gu+wnhOJGvR4B+yqLUjXa7ktuCiPDbMuUBPpHUbmKZJTN/YBYULjelCM6A1QvW
sZv6alJ+yHt6vVzjIAJaErREf3ltLRmrP6DAB+RD2817sQJueiPnPEu7UgnY14vZk1crBpknoQc6
yEZ6MNfqanac7XzfGTrib856KJ0iIuOjHd6YNCOCY26BzDYQR4X6jqM4M7OXligYXaKZF0S+gK6x
NONDmOipe9DlRLbyq9nvkQ6YCwUPxqePUm/AwHRw9lg+sByDSKeJjgi7saEBdGdxhDrZcEM87fCf
u8NNilzzHZJUs0bMRWffAqISj9bhc6N46xQ2vHKO9epxKGSsGhainOFp0Ydztkn0ujmVe82382Hv
xUL9cmZP8ibJWFPATqczeEsgU1nzMNka/NlrYaupQ8tYsKFuMky/G2OADvUJ8VbgXgFuakW4tlek
91MApbu0n8ztr/4XTjFibNmrKOSdNhwWmKo2UQXd1iUWIVuwxLYjBqUfxD1EAr3DgculIXmtQJth
NfjXVGPvn9BY0e1zunJMfaAhqJPXe5LzEBn9QdCpt/etn+1PW6SEtZRdjZGH9mf7mG8GeaMvEDMW
8g9GzXpQIAsESZeU3CENvFJSakeQo6rMH53wm7O9p1l9kj/AIEHOYxycI6sLH5geo+Qo+EcMeUwk
w7EY4KsrThIL1LgT7xPrKu0sSp4ZsuLfTNG1UZ7TCZcczbvZXtnZ3giwzD2DpBRZV1mozirjutLQ
05/3ol416HdYe3B9Eo6GBAG6eSKfUlut0cCKuIyCJ7qh+frB8P0j3LdK/PpU2G1qtbaipnxBkcfL
H1ajpB76tlbMMMZUyDnSqy0xrsTjudaAbk0+p5rf3NeBSAMQnTrIjlqU8cSrkxIJlXvVe+Q4SrRK
FTzdIIIprYujFAh0kjTElyFCnGQZwVBRGSMYSNAp/d2hRq6JVEG2d8xE39hyRsnHYdiWN87KjlW1
nMDarJsV9DtP/ZRxS8k2eQUKEtKqubiyCY+IOAK1P3HMun4BQaz5AxmQZPzWwYnHRJm9PnVm50gV
eOZvkDHkq5pDT+gStc0miocKzCC8QIDaKEEEX9kSIezZGH5o2iUTCPGnb3RDXl61UleoQeN3h3OY
j4ey224OBk3yrf+8JkktpfVegPPgMeb89Pmr3++lmovFu4fxvqsW5CueMWxz2831cTdjEqvEL/uG
LnUwAKLlGj1fYOQk5RTTqo9YGSOtEBFbxs2bsooB5b9DpKlf091OMhWIpL8FMkZQilTZMrczC9zZ
1MTO/pXtAHm7jcTBte/EGgPeEvipfnORgCnjqD1Mi33W6DG0MsBWZxtVIVy7LQrAMKY4iL6mbh1h
VkDC29F0ohpGP4N0VFdPBhVuymQA5VQMC6ye3LHwcjR/Z9oELzTL343lR4fCOTiDQ7znwsERCGrG
zOd20iSYUmvr/vIh7Jcshs3PB3/8dihJy+t/la5qViM53REU/JHP464k06JaF1GmcRtLUmE4qmXj
CoxtsovhVfgkmG7jXaxng8q8kG8QScnNRACmlAopG2N8b5VVOtc8Xx+/nqWPtABftK15b80+5QQY
aS0xn1rhsHTLvnjiz9BF+LcS9gwingZkb1P6SGIxBZw/caai4UxixkJ8Kf0Vij//6IN7RX/L9nsi
MV6GNI5gpdiydiGuqvdbL27J8yg6Qksxj3+Npl70G1ra+S9vCnMqiiLAszVZYLzY54qiJay5DgPW
Oh2mwwF/MdBKvhuAEJD6phZePEwnftnc6Dah/X5BNhJX35lPP/gZGSkh6Bkx9hIEYt2qIpAVOwE+
Sqxz2sZ4V+ONKiujVpeSaNvvl20A0OSN+29ZncZ0IeDnvYkJ/nry90lsMRijYWMT8RE4vWrE1yU8
N0Ham1WmQrO9Qh87rBQO+Mkwt1wcra4JNnELrfDAO/PdTnnN97Xu5N+gkdkW5WRBHyGpybr2YHa/
fF5O84FKVuhqk0JkTR0sQgVC6oayGhhi7tA2CQm1RZeehdnesS4Vj36fdaKtcdmITv+NuoS50s/o
VwNekUWVPiiLcen/NQri+3Y/o3B4iU/v8eL7pgoe+gxmwrHgnW7V2j66/Auk9SdLwSJ0nOfcSYPI
aBlVsfhD5YcbXRCwJSg4SgWVdjWhLb+nRU0+Cqvenq3hk1JlW5rpw1nAzd/uKpUOkU1lSqTeNAsd
JOK4iHbTRzlidZfYmHjW/0dItso8BINl+YtLgecVSIIbs442IG2Z0yvuaFMJrnCi2mF9qUckSOWe
ApGs+jsZDfmQUJkirdjmflfw0JuHNbTYZrMTztjGHV6DCnM1msI/VEgW3QfjNU3RFQ9XSE3MbOYx
OelPpkQ6nydOKMe9VucUzsSXefr3ons1NX05cye1tzr2rhmFys2VFIbmsJ+NwaNNl/zxsfrVzhex
mbCpdQ4TS1fxtrfD9fUa6h4FUX9/XORjHoOpc7vdZ+++2N282FvK/D6jSv/XT55YfIyGW7Ujd6mN
NsUSV7OejyTav09QQtUEbfGA6GZlsdVofRwR62jWdHqI16BWgVUEkGE8ng1zZh1kiVHQP6lSvYX8
bBq2y3PevuOrmuhHBoWC4cIUOfVeCCqs8MDkvxrMs2d38WPRbAiPjcBt3fXb+ABBfhyb2CLqyH9x
T8o9lUK+MT1hHFNQ7DUv3JXtK9uHXnrsP7cbeXszxYXXku2Z/ngYnWkF8orllntNXUmf3jk4ZMuz
m9e0TxcOWYbx2w/IoOSpfKC1P0c54F3y45fywDMLHfPijCFrEI41CRkdvs19PYorVsT4XECiKoP0
JpQEwT/ispdIr7Hkr2v2IduhGJdTN/kUvvO++Zhf5DNRIZtFdOvTeLWuDsa4LQTocSqDdbB/YkHV
6dlF4S1L/lcF6e6HShTWU4qlaqH8RGOrt+WLnlBTE3D3SMj4NfU1wZTwMIrw5G/VEuCPmvJ13VnE
UCqbKuXHBgbPcqu5RA3asf1Be/jDeVkaptRRmol1w1wthEj9PVk7gtR/tq8+ij622E5/ZXtSs7yo
yUNuD4T6URAnzWGsy0IifiS+buez9woIh9rXTS5KnDpfIwGtjR9hTzfBQ8b1P17+UhMbXhh8TOwl
TFGrn5Gc6neU2CnFUXuMDOMfuPBDTdCDG0BLcC0VzG0zXWAZwIr5rbXsSnxV+JTbN4lIv3p6JkRf
15ej49adEKldU4OIR2p4mUZNEc0iENXtVCIod8OO+SqJkw+gfDAZ8ZzOqBbRJQIfdhDjjUpPrJnu
gd05ImMYiXaxmTMSbWPT1Gh+8vjGU/gubq+3Jl+EHWTQbfG5ySB5N0Q2UENHr3uTHZU5DpQZnYJE
gLyiojOSIYJH2IP+FE3aGuqMhSMfhTBvAtYfTivXFrBgaEfRKnrLizKJhraUVufiLc1sKiDqXvtL
rYDP07LMigeMn6sV8p9EiiX24Zv8vGdBfAHb1y5fEaHffw0xiweJGZkVs/1pLrPCoQ20Ssa/hxkj
CQidrT/1eonmo2E0UGkYVPBT7L8dro7IxEM/+Vcvpz3qhl8b4oYq+KPmsQ0KaDTrVFw7oF8mkHVU
tclyeOFnDk1UGgim+P9BzbrhGXtvVFAfawElkBnPzHDy3lT6/6sT86IM5rPVwLzdCE6sahaUr94g
+cv0lwjdeVw4LpLodlj1fflKk0RxHVv1qoTnFXxVqsm86j678Q9bQjCRSP6dtempPtW4IBXosysb
Gbo+3TSxjlL+d0L0RIvHf9peXD+5MDpRvfc9uAWzpfFkF9KZjFv6V7O3U7b8weH1j18oRtDGl9FP
H+XQXOz8+ygayBr0xybDljE51e+Q59M6DA4K7XW5J+j2pRw0Xmnjbh1XsmzmPS2QaIoPgIIzkaCC
UlVT8UyW17TZog7igw9ISvGEkN3dD5ct354aLMTkEwZREYu9wMck7gryl5Jq3fmt9KpWqetJamf0
FiJH/avvDUc9rkIhW6zy6jtvms+UGAvCxtS3+1z2n9NuX0WJxZnFbMHeR/q9t2Peimy1imG7XvnO
98pRANQy9aVtaXAU6KN64+BliKFMbSb5PkdT0E8VkgLaGBOHLZPvFGcml4Bjlw6pxG/eaJI/2/6P
gMVKTdou7O7+gf/8666jXUZcN+xdZ2Uemp5UiLYoUMAJ5K+yYV99E75vvbLygISD0gc/gFQbnRGa
V1U0zw0Tka4D3pCie/yxqb4vV25cSaXau5DSIkQkcNPENhQxldDQtXlhqvC+cn1GzU+4sqzs9JyH
61p7qk8pJIAF2bj+XHZOMb6USGrrP3M5WYcDxr6d8I10QcdRLermA102LJHc8GJKl8eUTGxzG5SZ
oeXo0uKaKP4ukD3pdYxESWmZh5KCEuQF4NKAxmtt4XWSpF651ntEZLA5EECJEEoYe+scE7Cds/mT
DVSnvAKxm9Cdu5j3N/4PVx0YMnUoQlz7F5cgMLHNwL1V/vRHmSDezf7LGg7GQGaKXJYYk3SuJYW+
kxUO+Drgd2MF820GNpvjdEIKCLvHwO68adrNWE/RFPs0mEr6PkwH/fDDBhpAGFhfzBHYX4QDy3kO
XCw+srqMfIigYVMgzwvM22PRDv1pZAg92Ebik120O2y1eJ+NcxCjBgR3mVmhPatSMH3yNcwewOFb
BcWEitbGs9vNkVCyjd5AFz/iTXeRf/L37lm9OWNEIUiLhkkbSTlFRKcUf6FiBfAmu24u4x7oGdvO
ik4ckzT2/vl/RvAxprVgsJcGu7500cY9Fid3GnyRwdSAFIPO3vl7jHU0vuuKVAh7f/braTfIXH55
NjMJxhNXE/G35tc0K8hs9c9/ID6jewu5TJo9PA9ssIcZ7jxN3Xwi0qn87RwwM57PS//owEZk4E4P
74OV/wpwoIqvAPy2b10UfZLOpikxsY1qkh4hHENDo83wbxEGLcOA4vH7lmP6F2xPREcEZ6sX8mMC
+CDK63kq4ZtQbZSjBLJ1CeUkjOp78SZWAolkUhJSzDSr4QWGF3g9FLIfVBxotjG0B1aqzOv5j2xn
oNQEPDE1sxbWjYAkH4xL96j2QpX4xEf8gQHJmWnaMfMDPfxm4qSbeXpy/39vosujs86Vvs+hbLYX
DhRf0H2aC9Z5ew0/7hyeioYqUjya9b8mvcklEqXtnw5nIrMYD/bImRTmk9KkpshGLBLB5d14EtAi
FNYq3+hqGwPVo/PHbg4Fm7OqjHzoPXfwEPklzc3ATJD+i+FsB1+9KeONJq4D/ETTWYQB8tG8XiGg
r2VNiG6hCriXGbdcHZIsm2ptRJpxA6atvzp5S5qMZHvaUeYuS6Ai8DzajkYdkf8EEy8SflQAQnv/
hACzIe40ujEoU6p5Ip1f/UxT3VyHcnPNp48dsou03ebRvohBdtOekEPD0qV3n7KwyT7Q0XRlE1a5
PMRaM9LXCrjBwTUv4Np19/o2uBgm/9F4TqnNXi7bwJFZkNXoO39PD+CmPlbgtHD1FlFWT5Ura6zd
weCerDXDeJZLkuBlJZhyQdDq9DqhSor9uIkgMsVVJAftO4RXrmQHNmdtkk4/dEh0Eas8J3A68Faq
0k7BVy26uXPJTs/ZFqoljAxW1n0pbs1YKyRba9cKQAld+ln1N0n0wkt01nDI6UJPo1MUOaF98yZW
VA68CxmTgah4UkD6uD+XkfP4oqjU/WE4hTIn2ag5x5+ZHGbxRW7lErSbt1IHzAHb4qhXm753zpZm
pvkSiibxc6fAb3wkqmCeR9iIW0h8pq2ltArSxr8BxUTixcWRvWcXrem/Qew06NWDi45BPMuc6l2m
DOVhFcLzSXfDNfQlPfVrovRYoPqfGVxY5pcsh1DfgKV3NJ/ViQpIcHQC9AI38swUioY3pu2V3GXt
j20qNgC/TfeEol3upLvau9LEQiWdJwAu7xiGKfGtyVwaBRYXO01Znt5/BzL/KLzGJGAAWrVPRHXf
Gc5bbclvFiDkgHjhF2XtwLgnck1HKiXgB7wJkKKs1Lsu8afNCjpxGJcfkVgQv3/2fed5rqfxuAGc
4BBOigMM8m7WQx8HCoToAAnZFLARboLfvAY31wo0GQ4HUC1S0YPJnyjIvuRDI9bo397I2jvHsSsM
J6zZ3R/cbYlQottaia2bSWh3geFemO9ydLCUAOpSvm5T3jrDxFq4DV9LpndJ6AbYmK3lgxxMsiyk
06LjBf7YXgRfrsXFFyrQeEe6pB9TaccFBxGiCX9s2lyIW2Wm3Mr7b1nVkdb8Wz4UhvUprmhKHYc8
g/U3+KGjcCy4bD/DfkYOqI6itgaA5JyA+NBxEC1Ewd9Sqa4RW2XCNBDZBpH/aCr4r8qM+e2i5XPg
3Nd5SADE6foDtFRXFFGpegXYhSjmIg6b11B3/qZjO1UQJ/jie8XJiF66ndTiDIYxGAk4Bd3H2izm
wS7ko40L7lL6WXUJx/zpuGgvu2njONniGPL4dG+yJ+uOTzpJe6ymLokCCIYv3SX/n112QGMFkjSn
GNVMSzhRFOZ2Jlxu8LIs1V7hNnq7t7JCiwQzgX7LzWwC3UFhTNcbji1iL5kkMXEJDZgOPGmiYhz6
wz1LXWsAweCuD5dE5DDZLPC/Ry/UheGe4iQb6hHfj92ZBkW8B+zHvGqObAiXJ1GYOCjmt7wKRHA5
j6wF2XVwmR8uDzkrd0xMUhmyc7RNg3G7BW/7QgdjHVx3fOidb2V0cEP3nGyyx1l/5w9y8uWW5asU
Vw7pGQQhbEx1lxpvmMpFjOMhyB9fP7en7k596GWy/Pj9aAjfo5/iEEF6H21mSbbLF33SoPO8lDIY
AaXrPNZfSYAcdnQ3DELyPky2uoN8ppIi051moJC2xDLtru6PLB6C0sGbWfHmDeYsPa5I4g0dRxBe
WFORbN8ybUPUcypwSYc+33mKL+ztv5RBODTiURLPkbGw9GJY/s8e5WG9X3NYKwM7Mjho32OND3nb
J9dS5hVISZo1MbrruVjH3bNJf/qYKLQkHixUQQn6CqtGmx0VktBOCT7Cwd7rtTc6ApsIHGDC9ujL
aPH9mX31ngF0GOGPzOaQRehCKv4rPKVbWjgYNUv/FmMX5Wox1eGwBxehdORi3dR+hDA6CazPukJ2
Cn3otwTr2YwUXXy4qhiejRHdlAsD09n6Zg/t22R+vlA0hpY6q9vAa7u2exfcq1ZWVrEndqnlWqfN
RG5lK0fT7Y/i1b2e0vo586h8Yqhs2XHYjbc0GARG+m7zWP7WO3NVPgUM0DCzLq1A8leMZt/TYJBU
R/BGi+23IeV9HEKSYDnN9dq3PwwQckkffLGmQ2riaSTgFVXNCxd6EvHex8AVta+U41JlDCb4Efh3
z6yR3gfqS28p0yJxHalUKDbsHOJ4HofAc9ZQBwYAiOk+u2jYgTlg+g2ZRx/cZ3Yo7w/+PqnjTzXj
gLRQZTU7e0TAS0fgRwfP2m+dyByy7jrIk1I9/srVUS/pj3LW7V8m6hfPhzsc4huKvSKGVLRyEt99
v0Mqv2BZ4goa791THle93V4zaCsK9oL8oCZymxkb1r9UHsvKHjC4p5nd3VZxIeaVKnMs310fQV0N
ItFv6Z9W9/qQRwXAusTpluMQmMYD1RFrFYFyBA0kMW72y+4JVnivfQyWs7yo9Fy77Glw8IBZqyCA
Wcdgs4OlJpBDn8/JM2LaqEgBw1bzQ8eYqAHB+dzdgBUaB37c3yiGOOGjuz09pk1zL8zCCZGB4QRR
N5Qp730tEaN722kl/Dge+cpw0ojXlUx4TwrOEqBax3APXhJVZZwjLkDgpAqabKcWLkLG2fD14yKI
seEcf83H6swb7CgBeaWW46EMq8tbSn4fmKwGNv5o7Amh+ncbuXnl9vtQ6kAMzKsAHXSiElLLdibZ
W2ovF3ti1GJG1xyQ28xCMedC7NxgV468XtXkmD3xI6wmDcrRnPm821Ldjuz+HkOjb89QPT7+Ba/8
3meh57lMa1bnDxVB2nbhskIfyzxdr9HhmSNRO0QHBU8lRDfnPfr6Pi9ljom06QDu9dJ0eQ+NCm2D
D4EY8Yma9uI+i9WfA355xUR0uJOpPcJvw3k8tHlSXnatL8j9Vw82vl/jY0aTKb0dS5sZF/p/GTDt
pzmuQH1NcNJDg27LDa+Fags7cYF8l7RDaq0phOCbpFzPaEf0XKfYNmcoIaM+kkgPEQg27SAGcykV
gjYK/r3WXEXWQ90Ue46LBWmViCW1SdKDUX9TgfDvOyW+nz32rVAc7/V8F4NnKLvNBqJTgoWVTBkz
azu4iLsc7b0o3GM/bthtkinsBtqEgddHCzCJ66mY/xrABfgpFaCAquL5KoMpzhgVGYojmRAuWrYJ
gXBzcFRTVn5HogIMteZeVQaIe+dOyeSRgn6xwje9tTpYn07GzUQ+yk5QV2K+pKf1F4QLGeZMaKgi
kCPje1+BopbDUzmK2d+EWp/hPlx6hwFHzXzWYp2B0g3RYENwnjeA4WzWDHo9VM7QIs2QUfK3BkHj
c9z00UXL/rxr47PrDLe7Y9+KAcRwaWW4AroBf5p/fVCO4FFWx218eCRwJ9ylWP/9HinRRHzXgCFi
AFVbeGfIsfRJdOZuPazSiHlFG4hNnPOH/CLEOF/Ao1Bu+WLy7qq4uTOr7Nc463wBeg6ZDC8wGDz5
ROTEfULH69nOFxmNZKZz9bttQ5Is3IBrh5ccMjDKp0R66HnZVffYKGYpW3VD1eHwrxx+hl7Z5YwH
Q576QcE9CVCjdLtMTPj+4uehLXmNULOi/ivWGjQ1huwDqiwJRKzlSIUc/dAd1gve7QxGJ0gp1lrc
VDyHLj38MZE2NGSQyVVGODb7DXmoKS3gGr6cAhQxRwFGnNp0HBv0WrSsn5FRXXP4fdCylGkiDy64
ofj6ylZh1x2psammNSGqjzp6GFHcB/3rlQMy7TzSvSP6fiqIml5D2QzCnOySnBUqM3Eb6moG0rHs
XCsdwPkpfmhYzBOFQL5EwRGL9bybz2g4IKBV74BeE5Nvbtc9t44fj0q8xAYG3plfx1ZCsgnjj8GD
o0UU8eX+en7VyTy029Gk0GexeTdBlQInpgnX9oLrwyWBG1RrjG4utSWIANFHUSR6/epKp5U1phLV
F4wk4nbJ4tLOWcR0vW36Jwn1JaJFFnFjoJzGrV7ynP++VkgX5cRkJav8TR5ux1QhXeJljvY8GN78
1vVXQ9IqSfGl/3Z5NgMpqqCc+KGXvaebiHFexHZm5H+3bqT3HV8PGq89pPlfXR7tJzhvb/I68r2t
eqg2jpIs3P0ckbPC1rvi0fzfuV5Zmw3sqeBk7q1pyrF5ciKwqVGLNZczfE9Qkoov8hgXt9gg5HSO
Kb+qK/F1t2Sd6QdVd7WuQo7P9XkpUXokMxmAGfm3wREsTsosGWkAAk7md2Z1wU2XVHp9/J34Hyj6
AApHUC6y96XdXAmkKGkz08Zdktt5nP00hQcJ0cAKUlZL8yb+HYpyFgfpR5CMnZrtKj6sB0oCAmYQ
Wok/pNNAtAODOGJZUSQNWkU79nJIpq67WRFbIrE0Z3tVuo93aXjFknDXLx4p7mJCzqlNdwpDdnYs
g6beQp4aEnJu5PaEphs8Pc/ztUdMZ2zzT027YW1boMd2ebxCY2WwlyuX0OYulg8+jhibmZIWO4wX
63rZWDt/ovoPhDmi58nR5D/Ci9q8OcdflEfl02dKS+LYQa3BRqubxd9NgURu/l/HvW3elj2xttDp
HKALaOCKzG1B3COgGa09U4oJaDX8wsFWjx6POP6nnwY9vfbBrTd9dfObSssX27Y14aoBfQxGfqpt
OtKG8s+9u82ZXGjFsK1bJJuKBuVU4ucbZybRvBoxgwUux6rec8Nzgz0nW+rNYRJYI1MwF+w+9CJH
AL8nk1069PH7dfyJizDVmYFrlUqG4wkrLr0NALMOCAENbbBqs7KNCjiyJcVAePkG8TLnEXjbr3R8
vcxVHrl+fRPXuGr5mI2LUPcQ7+rAUZ6adGtpaLXMRpZfVnST7r3F2rNZ77wxeyzlyll1wotgSij3
zOPT5oQxPFk1i31iCaUyeUde2cCls+F1FNLGqhF43yUbBhgsHB/p0p11zj3DzJI8kCXyO9dNeKmH
X4w4ir6YCsI1EbwgkOo58vFSFkPVFKgJ9BoY1Qadvy3ALlma88FwJWuzVwWY9lWt6Oft9x4hFd9j
H4kbvySDXfczBIvVC5dv2+F3RnPYZj2r2p/LKGNcHn4Cqor1KT9lDhG+/jdtqMmon66ofW/+YYkQ
UTYM1tZ7UAWXvKv3F7FpyX+rSmpJp0q4OK5dr4Mi/cDeZHHxlRJzXsbGzk94oidC2hzvuLiThEps
CIEdXu2/kPmCZi414nrLPGzTvCjsOC6H0Z2riN/cMQkkjelfbgJ9Bt05k31u8OD3ouTDKjEUJPsZ
cwF1ccY+kQd/9YaqAMR5hHRK4QBiK31Fjqcdq72/OKdf2Mrec37KUfIJ45K9I9yMF8iz7O5T/Zrm
M6aon2bIjaMu7rM/6NbVmERdElmHOJ61+/OmjgAq+ptbq9kXInTxSNs9mifqewPFJqXoexia0TY8
ELmHxtfWnhqdK5hUQZc55/eaMCF8k6iBoR2aVVAlQEmW4Tu63CamgD+pvTUksdOM1FDS7vV4mv4W
okQEUJPK6LZLhe8r/H0KWZr2QnHGVAnXhLAHCuZ5ZiRHgwPjek0yslTY4yKuGF7XdaFN8IAy/GAS
dQYO4/rVpv0MsLzWP3uXZAX7lbCUcocXD3DegFu3jQz0428JLLxqInchaKLsmPQ080z9RYqN7q8Z
cHrw/Z9lIVC0tiY0FqT4USNtPNPaCUVuiZ8KZyOb/3P+aiknI51nPMftMlOc0ArxuBbR0KNvjyOn
UyPrKKK86xVLWVCW5jMtZudo5/p+zH9dBSSRUwH43xAqBQWMfHS0QrMTysaKWaHgbjZn8JGaLobh
9gbJX6WWzRjYvrXFP4icx0bBIiPcJntjz0h8f3/0mF6ysHslsZshm8IpxOSndFEnXmOUXLUzF/g1
mjngguqYQYsUU7dmBNj57qSLSvLQYGGcBQf42ZBJhGjZnmh2Hy4vyPtkzE+vIv7aSDlW/GBIZSoZ
eqYyxeq2sGaaULFCunZVirOLr7evRAw7637pwEltO/Mci5Q+4dpX/TRMGgtVkvipqOmFoXR4vBOJ
qkXP+fd0DPEseVB6SUKkznMmtViy1W4iP1S2+6ZpG+t2HOtYe+HFJeBU6Gkl/yth9KE1wtPuYSAe
9DtDVEl87gSxhwMSwaaZ/IMOEcalwd9A3Xe6Pj9zJbDmNI0tzl6tSshD60VOz0ZlRqXL4eO6bxRs
VBfjf+RNjNn8P5upplYg6bNjGKuKDtq5HiMjxsiEObOSAWMSlnVA8fMNHZFWml6FT+vR96cV0Nku
IBgdTQywWkfA9Ztp9CROXW4NV+uEdk33anlmD2wtsojYh+cmQVEsDn9pa0FBmtTfAHkhqkXUmEq2
xZ/RCuvxOTPFoiY0URGLYRztj2DT/RP1+Xbmg6f5Y307gqdm2aLeDO2q4zmfozOFLkZvtvr6MD00
6pAwaEw88/c82EAENosPCPsx4RBhpo6VwYRToGkcZcWh7x/QdYcduLXrYqR3s/VWDiKRxNWto4+c
4O0SR33UUvm25FtKa0NmFLiT35HBNY5HAgPCnIdlIPE/PcU+WPhx40Kg+yKcyPAQM7oj3LohQhU5
EnQH83Hczft+cCm8x3qg4ekvBFhrM/Ew56/ZFSCYXf4yX2SvOjtbGULLvu84VtIDT1PyreqMTYkH
u4TErlH3sZVrV01AiRq2tS51W5jhl4MFq6weeUXawaAHQznfOllLK+iXF6knx0KOZaGSngmqZPhM
db1CsV6ZTrjumjhkoMs0ZhM8WrKGzW+9JRrXoy0yckHxbOg5HLDBWAFSWd4Tl4waETmPx/QytCiv
+9FT/VGXSSPUfSbw092jdSgzQf3tGB3OowBbEfFmX36zW9LrTcpkuEW0N98gYiOSuWywtAVaFAwq
lBtpOMDPhp6EHEmssIr4rPTPk9hniO4qD7Gw979HFon1q8XWEJGMo2r/YyRwrcQUvIDGN3FapXai
7rvpEarPcdSwXAiBP4H//BYLGROg5jr8fyqAQX4j1GtiS1yP2Pv/ceK7I6vCukLzNH8vrEUoFxaB
6xjXr1RyVv8s9k4YSXYPnaWZtTz/TPVaXY6AF6Dt8mhkUxPxSwMeOgDCaSM2Q/Gp9ThGVXYAJYGu
tbdL8Qu6TZJmjoTPb5s8O14K/C4MC7gul1UpDI2sF6rHfVB/qtMw+X/kN717K8c4L0mBJqSoA58r
6ykQrFiylW4OoFJo7lZggER414vPchpEfinCCIS5f0DYY9606XL7TRYMuZJmJ/bxoAT1/1zuFIRb
FSiZ7St4ekPnWthBc5QxOplNqk0weZ/mo1RtyOQDQhkHGKqg98k0xbdeL8Tm8VDJKIrm37CcP+bA
u1xDnCczgIdu6BO9hC3kN3jzxrP2W687GzDFm0mOf4/P3a7NodL5uDjYf18SozrbC3ehd1GHZuKd
d1Remvw+usA1nd9yZUQ2Cshv5VS6ScWHsvYT4hPLfiW7E1xPewt50RSd0JXfJHaAuQqdfxkN9/0+
1d5BRHykI1e67OTJGDrjMj0wnj8JDNRtuubcGGYTC/fDPulifZLVQIe2pgFN+PnhZaX9xSZjMANX
6NOpo7UPFAcg/L0p4b2FbdeErmTr7WQ1YPcwZcCMo1ZXSq3vsokvq0HRXYHqNc14P4TVnHtsICwX
7o8lPhIPSBdZ1GW4yghOUK2OjgVcNkbT5AKJLloC0LxbIOs82n1qXHvOKdRelSe8CEqtrDGSmY6y
fvBsR7ePyaWK2jewH9recySzZGJqUpCPhCJF6xk2ir6ku0TxDaqWzKPRDUOBJeV1N2t6F2F+C+O3
j23g5eklJEJFMATcQwW0Q+ysv+iZA6vz2pwi448iuaSoJ6LTi36t6tHJ+8eCUpCO8gnpMqceGRS1
aZBJEE+ZG1gmcI7pmxu6zKndjfaLQqHOmsoOprOCiabWq+QYTFeM09dCuNzcXyH9x1s25PjVywfe
+rBoJ2iySP3NjK5vHVDspc9DJgSsqvOoec48l5sUelpR4GJ79AFQr0kugz8kB4GRIQfggg8hguH5
7zzs8O0QOV+lETDUzjsvZU0aWi3aQOz9INdomv51SvN2hNMIBarBSu1HGs/xOMzOAbNrkVPbxo1R
Oi80z+0WV/MyQomL8ShQzR7dir467nVhIwBfhMjuAUhnlR+igJN7JsOVRCpAIMuodcCfxXroxDev
2sgK/+4PR4R4vfe5OJjIXp82NOmltuWAvNsQZX4j50LecUyl78N8QreyyohcGR1VXrna20lyX2B8
GzczZOq07huSmyXVldbQHftEMPrTBEVnbZQu5Kdy/xVXdZxTzTLS2MxtWkaFal6A8TnGAm6s144R
L0HaOIdKxOhJ7Ux2WUZbDRZhECRdILKvQxfCOE5yoU6p44cYA3DZQW03lPByMcA10ct4vHLZqZZt
F/3CXdLVNMSMz0U8pHhxmeN7XZc4ogylno4LJZXmbDLbNewRN6hCtIoSUoLq6G3ld1QxXLnBp1C+
6Ao5I9BQ4UmOpYZfUftllQeo4ClDrZqFtfAckKINgopyIYfltbF11LUWMe5vSv7gIbRRZSZL5x4I
EUsSbuOL+WyInFFhABu0A2tT+a74LqWUrQS3DV07uVbZwEAc6sMqA588NHKDNM/Ie0QM/wh8+pyh
/dVhjBb3GUhCoKO2PGI70vpau21GKdm0q/F8+AZv91OvlL8OfjexGcOvvGdmNf7UhzDVdKjTckd0
4GDOeEHRrG2HGjM3isOG+Jmb7/bEQio+oQLx62pv48g3IOpZSEZhEBlIXIN4HeQwnlKmzqdbbEnn
ogMe0TwwB9AsZYucEGI0K/woQf2+M7OgMad26tKlmw6IiyX9ikHo+rrl0Qom4IQuH06AhwkHseqv
bzxZC8ScCKOoZEhnS8WCB7l5/X5otW2yGgzLh1WaRDNi0EXpTmB5Ru7VjIDVrOoQMFiugKmYWbWg
+4Y3p8pkS6G9GneLriqlODuP4HzP6ItuO7tlAis8oDP6YX2FgnyV4Xj/dcvLp/1j5dyICgNGqSyn
//zox1ZZZd4ZAsryImmJaR055sdVJ8x1Ne9Hm+lq0+AiBB+Gaa/xIJbq2YZ3rBb4t1RqMSGbz7DU
CfcQAjHnmTCngVA31K+lg86nucP1roH6oIAJ2Dh49daMw7iaNMBF3Mox2kRdc1ir4I3EvHwRRWdp
i+mjbctgqucgNmoyk32b7JO6zTPnqxt153SzI+5Ndn6Vc4ee4CO8VptkobYFkDknSKV7nrQfPhLC
KtfozS0HouwW/crogVk268v/zoYw9ubTtY3BIdNAnqecuZ6aiMfZgdpDme3Z7ORt3WdfIvikLt39
aSsPMaBfbTz6oFOzM2CNDhUhVkBLiMYr8Ok6ZXdMcwR05RNKw2NLj9nJZ37U4k9ANyE2kVkqYX5s
3I4LC2SI/CC0IS1IspyE/JVCib1GXZacd02fpjBSJL2H101EzwoQ4hivVk4Lsfwm7OssRJMHXX4x
SvBxdAGu1VJQ3E4P5IS3QgOSjiAA8WIaMA7ZCURNnrt4fdMyHrLvy0W0+t0PtgxpYPFKK0p3UcOC
xHEM2ufCgg13dBV0BydMolbgF9owJmw+XWIho72zhHMvOmErhMC7hwqgn2CFoZl8nZJCE5QUw9na
2eR/sNbYFiKOzd1bABCDj+z8IkasLeE0o1oA3NdWYgrlWnJkfvOHCIbSCAkLmjgbX1MltZbcTw19
rCCh/Zd1quGF9Kx545loLl5LE0DxawWl8yKw4PrYAC5QtULdY/1/M/V2CwgVnZypd7Vyjg+cQT+J
v+Ci9bKdBMLV4wwEblsbyfia/W99u/00AJ36ThU5GG19DQTL9pkxjqNuyRlEDBb7x+NjK3u71lX5
P0x9J/oqGZTmzpBI8Wkvc6ZMQ3JbKl/dp9EOo0nd3MOICZ8XcO2gqfnJgOZc1fMhjomzW2Mp+4vp
9Nu5dnuv4PaDzHobG650hVSE8Oq1BmDQMnrPTKf2Z9UKFAgaXY9pFJvDZ8OM4yxY/I3HQvVbGYmm
OZWMkSs4Fnk0Tdnkhwpxmqjyb6y3K/CjBVujAue+h257jH19zFwGSSE2xiO3YiyS7Y0hO53xEvLi
NfIxd93gsr6J7SkeShI6743Do4O/BLddLz/sAPq673XzPF7nZbmUTY58z+xFMA5FQHYpOOePO23z
fJgXZAzTvWUeTdQ908yt/utUkYxd4bBxIyAmkiQUCC8azvX2ljLkVdsPh/vESaNMvYeCPrZ1kN+2
a0+c0RUUy8x70CJyKiIMzCVReaiSyR7er6SEU72kWE66xe/9Ue9sVWv/espYyljZ2RXs/WxZJyzy
bTH1dJan4WY+VvJdPlCqyrZuzQ/Lk9+0gN5qWmnKbSEi8Cbcwk7QENXV68UQfr4KWz1qclsKvc4x
hGn3ZzcLyihld05YxqMvSncyHg+vn9FKuiHWcz0iYsXMpvz9n3mFmtu9Ve6mdb9ULkaHmgyHCBw/
WLMtl15qqCnY4kpmcQxV7860i5myShl+pHWc+YaVtkMUm4hbZziXQafndmjziC/+s39rCir1MZlB
qWoFsiH/it7HFoXpvcGzX1+lz8cBh1xCehFItcw4g9uUg4J+dWG4UMvH8n/ZEuvqD/4y9KC1i8DT
tEckOlHyKvbcm+gKt/vKWj4VY6ULl8PwDjXaFEVSzy+PPK4EO/QLTeJF8/0rS2eRpEC8SCQKkhwR
aZjPXz+8NnGAn7ctLEkmY3M8S4y2xUWxJ1zNfoATXiICa6E0Rdq43cBV7xArtbFCD0c8mcuargkr
9gG0v9uPCqdhEBkflyRLhn02zbIk+pm0BLeZfXJyoWDUVgEMG/yWQdhIr1TlG48inUgtcNHlZyyf
7sZJauhczqobkr4E4szFIXdO17TwuX5VNoTDwplDlTMyiQW7VZqAUs++MDbUaVspevgGE3ET0I4i
Q97FYacfb1lLMACRX84awy4iMM1h9e89TjHadgPt52F/6LQJeT1MYNiO4iKEVnQxrO4MdtsXJCWz
CU+hcVhBKaDEV+wN5Tr+/iVuaOY/ZUzXcTuHq5nBEgFzfCxaJldmnM2WeUncJf5shETthq2r7y4U
hSwTOh+MxZqIeVL9iAcBObAwGdC73IlrOgIYr7u4dm+6VJ3rZlebDojAp1rp05ushTxFIYL7xq5d
lWazpH7UEvipPdUiaDlW97QvZspmlnjN5E7OdzccslbFnFx1WYIpM7xC9OcjNg7ChlmmAPMD/CI5
AWrtUuIqWDSv1zlw3d12YM9x8m3x7RilSCsoVd/t1WIxROaGjgWjK69LCj5p3PPDTOWMi6PbVBvT
7R6jtwxuC3yLYFBDMMOyJwwovCuxceEk4LFjt48wRrX8TMuafkvGV6M31XKpoFhepzYjJ11XRiJl
5gPDzoTTJLYBvZ4Fvv3XT4mjIakMm9neJboAo2Z2uHIVDOjcQfYqMalPd7NjBc+hzSkkoESdFSdW
6Pjn41nI3PRqHtiDMEziQU9ZvM6yva4uQJ+uxCRMrPlJ0kMkJjwqm5PUgMP74Bx6JYXfAWfP8BXG
JNfrmMhqsxNubTfvbLcO4e8LFTZsAwCb4f/AUr0vleUZ0o0mOsB0Qy4GZ+cfOrVl9eUIq+uCZRfD
DwGsuDKKOeeZT7m2iJz3c8fxifDMIFYEZPMIRKIyDEtr8sMmv80HVJmoYoubPgLXLyBbU3WH6fr+
POoLl/j6SUgYfI5IOyeQw2R7Tv/XBgfKlR5pu29fAJqz1eXvKkekJluCimHvlz7j0VFsTTTgjNuP
jgSs1u555oeu6OZfwvukJTrHDBw9q3GC8WgQLBT5kyGEyw6MQlt/g2PMvMwZWwP/S0INPjJQaUFR
dg5hpOTXNc1xu0x6UbfJ0ftkz8E1RHfyPomoFvnf3C0Ao6DDjLLvsaxQyjgoNo/K9reesDCqZGIv
TdPY1lXZzyDDVrMse46JoaCV5yVSMzmlOu/90Z5Gb46UJvtnVUFlEy9vrZ22mhCGd/f4pT2qeHVT
KNgxSPx/aZJ+8bb0oyRcFbKxUyOFB0nXPM2oqCcpRJjmsy8vv3n0Kr9mMJfLtcprDqMDl/BcMJLb
y42aRxVR7bsEFrEYB96EsspbID7ZZ96kFZGKexmqZvF90MQokfUqcYb1BYiTADyyZFwGfrJkm9ox
w1Ght9A98YqpaE5OMmk7xVRWzX2FU4BSFFqZKJGPFVsPLnBu8T7ZlfsAeCPAvI1CQ/0I9m5ZkFgm
hVb5jsWS7HZO2FWvNzv5cUTU+1RJW98Wl4xArcPylD7pL5RD3E5zjLH5sUhIzFPoATgYrxzUnaeF
7cVravMsstFbt5O8/P0FV+0tGuBP3QqHLQ012OiNSTY5QJ+NNsgq25FFuHMIyQtbwx2eZ4wQkWvz
trqnseZvlpGvmDV/a/fdUnbHT1SOfN4OL7tLL4vsjqCpBwpa2FQZIUEV8nvw43IbQdHMvF9V3ThO
xPy5guBOH4mWC3x1QsiMWtb6B+geK4dlZfe/wV55aLlsd0/KC0hSFvDFVt0ZQUYRgqr7xWrZhwBS
YoSf8xAv3InxBkX9nObDklwLOUhqPQxdSmC+6ZqEznQnyh1jeyYvZWS6sxofHYB/k5ApWh3+UwUZ
pliOLFBk5CFLWq7YUw039dvWGBtyhMsThhqFHhtvxpo4/Y5oyvS9dHa9HtFzLFXH7Ze7VGkerFbn
LUku2Qix8smWxSdcvKtU8eQu6616HO6bkx7OqIEM+F2+HgteXkwA/zw7exy+0cH0GzVWXfTSzB+6
mQC8lnT4ZuKLrhH+uLe0GAZE1VDyRBsnT8FbLECqRPC3O5W3P+KtEuZ87k9stP+aZknkIa9yedWn
Va4dpMbhOg+RWD3nre95UBitjZm4+p08G3hwpR/4QZ2EHrIC9JklsJ4Ls4de3P1gGVf1u6r5JOVu
DgJAoPllt7H0HccNzrQLABCySHbjm1CSB+bmiFSalOi7xPrmpROKwYf1gE4D4KEyPhHw1QYITViU
gypW+ohvvRDDWxDCz6618+f6m81VjMXTJDq4aoURBHY6yZsjwnQuGTq0NALURExuMz3uygDnBdzU
4p9xFm5jGLhkdtlNPLqqQCApFiBuiYXr3wgCjJiZpAkqoM2vUZXGzdIKrVB8VwzY76a7+xFgB0rG
3EiXQZNSQMyQLce5zRLgYn89pOjeqjfeRqoQQHE4yd8GnWjNVvfmVWutOEMtSQtlgvRmuS7Q+vLj
cJZVVVFojnkB1p72R+1PE5Ki32cW+pGdRFsgIokxGyx1GQC04jj5p1WEiFvsnzlb5P/WGO4qFJ7B
r4JslirKpmSTuoCaIPrsSnlCjJIyzmkb/aSizXtO/7KgL2hM4oqFp+iv1+Vqnjay/h96qWZ7e4su
rP9/47DmdbjBDyfrvaxZYE6O9A87FxL0uPhpxAOfRGQ/+yrkBWyOGVXkKqxyWyWBFeb/vCRIuQeI
3R6FtOVhEHEe153tHVw+fhlSzHPeeVC0pnpVN2vJ/qivynUvWG9QJ/I7ZFuCkbZG1AYcDF3p5cnU
Ulq26s4nEf8z8VB4xTlUzZdODEcTyzWXHUheiC5BoBIYkuq2MNlYYD3SGy3Z7KmdQrrrPZPmM3z6
8hv5Mz/SARnWK0r2zMsiYJn0Q7cXXXtJWgR926Yhzc7kkf7jV1Tk5p7p/sayh0WCEmBCN7vMFjtO
WQk3QCbPysocR1ygskQbu7OZfTfR3AZnEqndHpTHkbvo+Tgg4nlgZNyI4S56fMNF6rZsAe5A/H+5
Cj6rR31BBbhTENK3gJPydUJN/Wh3Wo8k2WsDmE9AjwCHyS8OttDrMJkmF9uH1yLTozUCF/CKF3V3
E/SxRpSyr3PtA2rHZk+Ko6Ie13k9Aj/e6I/zSblZmNUvzgnsPBZv5jEiM1bNUWj733ecKaP5cI/v
NAyUlZfS9oRm+zvcB2J6sjgT1GdwTs6/VpJSbtBLbrm9/GNJ+PNjVYKzK8MpUl3VQjO07AWprw/u
UleIg2XU6a5al69izI7Iko5Rrr/APTlJt8JyWTlUps5vHDmkt9DXrzBuOn6ACTtrC349ANfBXtBu
0s015S4zdtqWxqZSHfs5jgvzNcHyL2twdtmxFWgOHRPESeC8aiiCYHxAlOCOQr0FwaxJcxYtqmro
SVrbNrKDdoao+L+3aqtsMEX1N8gK/WNewBlAgVx2YahqKG5BwfWGiANMV2Oh/CRDAv2fm5yNmfbA
jklFNfPHULe+MTUgVGngEY0BP8X9zlRpcOKQlaZLjoJEuBitu1GrzxZ2iKAUCl2BkTs5LcH2Py5H
/32xMD94qSUExIJFnhy9kQwdEbgJE59GZLcLuwRb9e1UEJk6n79B6fgjnFAKp4MvyzciLfrk7sIN
cqkM3jyV14ViXUAz82vA4Hs+dDycwK1cW7+52SKyJdklccK0BPl48ar0j1dh/MfBFEzWaS7F45rv
xvEPV5G4mgbN5IyDg+Elog0rsgdahNOAbZQe9JrZ2uXvAirpxQaNMwsxa5VLkUwQUb//XA99kjLN
j4jZka9eScfaR9OPbIw/3rxCzDVGh+qQyisJcMX2xqV81sy20v9LeXP9n2lYHVeMzYSsbh8Dwl1I
MNADO3At3uKD+T3BXMBx2XJoZmI/xGsasC0k5SBj4tBTN0L8nmHfSaREsgnOFesy2tVlGVigAZE/
++6i8jigNeHSL2BX1qRdBKid6A7mJQfujB50uDFGLCMNqrEoDptljqw6PSxwPBkCva1XeJtfCzUj
jd5zQWjw8VLFGXAI5+hQiCjgDdIk8klMNswe7uFFTRuYHPgWDFc+mCR5jYjxovMf/9m3em911m7a
3HPybunCdV5fhcm9Yxk9JoGidHChvcjVRUAEuUFHWg7QfNfXFMn0zMHdrokqZtZoESMtkTxWKxXC
OD9NyBzDzJG1WssKpCfzevlWIlZ9mjSrkh9qwOm78veVRkn7XMD8oImhN3zlS++8VladlHbF3ni5
b+KnNDVKURkjimub+ePFpP3gizrL27/Q3mN5v3uATYrxXNdfn+BoYI8mNpjG/JLheEx/CTSIiKMk
2sOfh1vAFdvl1kA9N70u7inONvm+C+dtq2/slBrpxk9mkoyJSwpyrcmgXQpQmbXPToy+yO8oo6et
m1m2y4HfZJMUQTpkY6v4FDffqkyRnSjoqVcLZDI7MBOkYPb2cJXKl5c6QOhpyF79Vk8RB2zE0wbl
eZgFj8jX3k9V7gP7TtukC+u0NCFCHkTjsx5th+DJ1LVMitzhnn7pMvtMvLGCcE+bTPTqNQshXLh6
LD6xL1QRHlOK68uFjrES6IJ3erkRlQaLPT9Cfpjb/YZ3nC/yZKuEjW7Sz6QvYb6NQKVehJZRu1Tx
mdqHrzo2prwAqaObdoZvZlb4ew+nlZX21885l3aX58cBlxWIf2bdCzwXKpq/OWaQC/uXtF2+iMD5
RViWd/c6owIVTi+3anOUWf2RXqsCx/zpu7iy2YLKJNjyBneZfWvm+GjTirbkmNv7KmLy5ZZzJglV
E3hLdihlCi7R3z293NKOzR6dhwwkkCSrusZOWO1IB8yxBDBWEBRqa83mVsQug/g8LafeWrIv/VJf
KzSyhVx93mH1q4yLJxwQc3Am18Oj82SVHPtsEErJs4tS2uhrT8oxwEC2Hr6Ng8EN45V0IKFzZl/I
ndP4o/PJPuZ4cUhlkIuyxi9POYuXIEvubeSKS1vgG7CF2O0cKsSWu6GjajdPab7p/iSLU5R1tTKY
ifpPUBsHWhmofPrl8iKAFk0GF9LsmdDSI8NgVWDCQMQMPFzzpqBcxeez6jbdgAWbWsvlFL8YyA9i
4peXj5BE7I1j/1JyTmW49GdGzDSoXcAdDExNv92Fhha0w9+ORhZRugzQAsioJNOQtWqGky2A7UQ5
NDLOFxnUon7xpaXSA7Wk7WtU0G9WR96F87ihyQZGFIPYM/KN1x+6bG3XdsnczmibntKN5vM3npCN
kg0qdxvQ8Hqet+I7PnyG6tsHvKDq5nrWQeyAk6QudAuMrAyZxptpwgTuYupJgA+AKaJAGNeo2Fjd
QZ+Ex7HhwH7NHSeBducIdHmgo4fkM97RsZ7M6KvUcBYN7/pDaG0ckQGCUF+J4zeZF6AP1vee74U6
cmWOfclFnwkEsVPnM5I5giGNC8Q4z0PA7VNaryuQfR8dPyuxH7I5m1ebJJcG8DqG81p3VT94GvIS
/fIArQ4QdmXa69Qi7/dQtopT7S8B8ZPLI3CuYqkizSvhsF0SvjsdYI/FksCfyawJpLIs+MWWo5OU
RavykjOkE3nHWheJSebwNfU6eoqVguMrTenCMNmRgekMENLTeNVx4vtoW8DsSD57e2vDxzLNeuS8
cZRqBvuiNg0tFY2sW9bCX9levWrAT19iDokk0sodFhwj7pXh515c+5fjRyU9jYWcVBlMKA1MPPRU
XQZmSDwtCMkjDnzgp706XlPWmJNwYcWwL2Pjufw6m9A9mlzubFimuHjVjPgwovvxHtqBng4otrpG
hDyIfdARmEZL3wkApsbc8ADf6HYft7iW+4q6aUb5wJKVsf044j2K4PXpF6b9iW1otRU/BFXYEigo
wrDSkl5ZbrSDdm3fEhgRuyvK+2fkWPBXQKJOGQ3Z2tIbK+fzV1ssTEOshu1KJaknM92biITMoZZQ
9vV5KnbqGQEM99v5QQplKh5R+gDQ48VmIjb/Lvwjr3pA4wilVsQzvugA0iD6+eHvL4AoL5zP0h6G
C8skV/3ipA/UAgVQ8I+PwGqoWPDSLzNd5TV2SAu6pm7E7vXdqNwr5eTAukythOg4w7hVC3cRfATi
AxQ96yTgaGxpF9mXz82X8ZIrjfpFIyWvRwn1JWjhZaePCqcSllWSzMOcY4WDnRutxCY7vHQvSV7j
wg8/MWN+dOG3WPEcjOSa3yNGLt5feBXfTZDtm6yg/vjvUzy3ykzlhM+U+7pWm9PQflbkj62r9q8+
SJFQmXr45lwxFu31RnqcJLA9W3ceyaU2MMzWG/CdwtxUnsEbUbyYthYzMvn0OcEGlqGfye6xneRT
nCho6O+7gjAY6wrJkc9gi6Vghqx2NElZpwxPATux2FTWZZLd5fEBz8Ov5HlO6JzuOYo9omSLnmaz
pDCkTmyfWuIXfTLkO1Y2FWigwQcntkUixR0y7B2kZO2AgZ6AKspVQu/o/ZfjP+wEb9M5y7RpAm79
4j0w0FRVBa3UHxkIkMcT4ch/suQxZMg5lXcPTko6LFtufpFEq5oQcK5jry8SWS7KU84wirZRvQK9
EE1uLjH0U8yPmgWv3P9KyOLtSskYGjDzgIWF8pbX+xE1X+srap9UdseU6TkW5mmj42G9gyYWquOn
g5GWoCoYsuRxC0S5NuEXqM2PtLV9pbygPnzR/A6pvBTysrYzWnyGXys0zl2P2dLaVYP60x9msRFr
mvumfaDasINQjC/EsJSMIYrAkyCdZ5SRcoH1/MxL238M8cBrAqUWz7c4F32jG5FcNKlTAW6W8AYH
juP9lo3nTSCUgd57BwQr1mthu/9l07pmAXKXyv8ipZS1COh2UrEKkTxdTQWJDTKMF1fJbI2NAd+I
cRfUCcUn9EzefegmIjO5bIIt2bMvOKEHJHBBsyp5BpLTA0xZ7DBkztfXSt8dHq57yqPr6K6ouLp/
f086hZ5OLuT25kJomgAb2v9yHt+p4C1FxtnABAbSmd+UAubxIbwbY/L0mHMW0vhXgHCnYwn4juPO
0CZHzCLaBWA5VxxH23jiMhnBN5pfOVOfY/fR9n8aackAcJyWwCc9XdpGyulb2tmmRNyvAvWhsfb0
bF9VUQ3Ijpfak/2IRbxgtOCElYUV7BVld+9F+T3vROnSn09GyAFJwiy/b4tDH5K/Es9iTGoYB/fa
R2AcMgiidSexHaQh1I4A524UoZCVSiwothUmHRtPRcayQNB7pWI+TLGsxnVWKLMb6WdT5pq7nXiL
68PkZvcBosWJGPzIBEKEgexSwIwH5x2Gc60ixdnr5Rkd7mRzoqBLsUWYXkPkZVC/8kfgqbYyx/Sq
7ZZb503ynfxl4hTWcE6awytj4mW9a/suoLEcp/2l0KhTPHGtkLEnEmxEQTdafGuQ9FGnAJiu3Sgu
MZCT865bFVzTFksz4CgE3NDNUm5EV7uvMlYp8XBEM7tNvP6wOB7olcvXiRO6XPlrDkpubhVo8PkP
PkEiGlD0UZt/xDHfSXAKDasYiqvHLXRkX3OTpZXHM3OO3V4srptx3itTFUANFowCI3nTUGeiyJkl
4i2/LyvjH0/qr6Z/bHP5fbd0AtOl7qsiKvB3QcSKVtztq7bFaLUbSBt5Xbqd7anAo0m8rVtRKCzx
agoM7NoHkg9mFnFRn1Poo3i58KBO/BnsYUc5RvLqzKEcnfpuxUYOpQt+n3/7vG175fxXzVtQUSBK
YH+QUrv88vKtppilYYmJuD+IjEsMShTSscOUE7NKVhMnE6xoQA3zHuGqurbgg8Rna7M3VYwVXzaY
q0gYL1Pz0+0TpvJ5zYvFdDd96xoS+z4MWayOYMmuQQUwhs6ryLoXNdmPx5EMFnmqwftfV9k5E8GH
JpTbkYLtNuYWRUpVCpLBHOOTju/GC/lZa/IcJOLs44SG0K7ZgaX09l4xDScCG+kLx3jv1FbsTMCe
bWhcbtOTzlzM1uaDKmoxQ4JN8R0MSJQUOAbXEtOPmuGhhwfaHh1y7/Hz2IRj7mL1RNkV/I4BMpH0
tD/OIpQEiyfrmpgfARAMvKOcz3OuXrVytXOC14vk+qVdzpSBmYhT6k03DN/El8ZuebACc8bgEFWx
Uh9lbAriGvWjDB8pZ/C5I1Ojde6SVLuRnwagSpLLSuVrp+LZQm6rlhtvtfIz+92KNi0bYuFkse2c
5z46ryglZa4BodOJwenyA+pkTRar44nK6WsP7pf1Nya9bl5iJcNwc4zdGwaNW6G5iBb7OaWP3Pjq
xp6yKL+gfGCmBorUKkv+jNwHFqKx+lUcuMvOskg2C7ufMu/WAcOnz5eB/Jf4d3gu3CR1jRiU7r4/
34LIiZs0SQ5S6US+eNhETJVeGbc2pnHHI/vsn6NwYlmBbf87uNcxCCjSR195xg1yYkR4fvMIrcuB
5EM5qQzLlRWf37v2OH6DbQPxFSqPHroLBdLfOEThVmYIqOR26bL3Fc/52zmZo+KpyXlHWiWCxMdH
0FsYUdufejBPP5pebhHsfA5IWJYgvCzBBJhxn09mRJKqtiyUgnOJkLiqQMcJqgLoAvBoY38V3MuJ
VHuXZ7lws2NRZb44Di6Y2eis/Otzl7bkENoeAV93RtaHYF3042ftaTZ2n4UzCP2B2ZCiDwJi4Qgr
vNWANx0qMjs/nhnMwY4qXtnKLxMgNo53oZUqQMDXwjMof0tyBNJhlxcYiy3DfNKV0aEV7zym4ewd
jDuxE1PJub63Ue3gQZIamVXIadA3oKieOYob4x2JWxNNriKdHI+VtozSzboRrFedovuF0EPZIamy
MFEV93Y01oMDBEEHPUUkmxybB7xOLNyUw09+rOZJ9Do0R8dSYt5Ggqzietj7vDs3tUi2N61X9U3n
qfC81xJ3f4RlNkAc2yqywdTBSpyezpBEgIiG2BiTO+CKSdLQa7qp6BtSP2EVkmKehxOFrVRsavsg
SuXNg3WuTeWhpPaqs8iEu7Vibr5KoH+9a0jf7SOj3tWHEAognwUD5pvib2URJNfV0QJlrz5y7MuG
izw6iUR18C1XPiOIU/HyqcF8blmbDoJDbM6eMm49TOa/wzK+qokrQCuQBdynFcSvdfOhMPlYCFuJ
Biap3cPwpus5QSmAk6fCohvMS1DcB+A+83hYwgV2dqZoGBLDErsvW9LH/V8GrqBNy69XpiCYTVLZ
yuz4EmDOTK2Y4RUCEh90h9Urtri9yBRC+nRkT4zQAjrmsZyLd/Ecp6I8+xiQWmg1gJZTbxZv/Teo
vZc4fDlxAuyekcmxK2effST4V24llUZtBD43Q/4Z8GC7lc99SPK/9kVTGdsfl7X/YBGWmlb/w90e
CSiUXWrQiZzKfdzZ2VNlgaUTu2fOObSEbbf+HMqBu6ptRYThrlQO8ppqicz7v3fg962/eQJ4TRSZ
NnvqUo1vJPE/TNh2IJwW+t5J6y4eFA/b6y5NrD3r1K8tE9mZSMB/inwa0Z2WfcVMrpgLxDjWVZR+
lNy3/hNCgjj+BX1StDQaxbM9YAokpKN2Jhs9jpdHCoQ2qx3k3VXDJcgkH6VMx7AegJ5+WY/7YxVv
mlJZrl4yvY4qnzhfXif5iQdylML6grSVz5MTT3VktPerWQaVAbQnATS5n0r6o8tCtZbhxCV4J1WF
Z8SNpSQAovH4/zfFioIYUtQubt2pvYGynWbI72Fx6YROJ7N6A/cU8oDd+IV6GKMcdcJ+5/Ionoh4
hxlfB9HdJvBVCn3mwXcG4eLsf+6+iuW1kYQmC2LcUEH0YPBR9y9ESUAJcVCmsgkuujAhhDHHULFW
dL1Dp21AVtO8h9bi4eyinrHnJ4HUqEf0pZUyJZc+GWRPHOZ02PPHCLV3jYqaVaqijNYgle9lKBSo
0W5HL8iFlSIPRg7Ms7vjgHtwPX0Wv7B7uHdkIqDcbZXGNKIUqi3Njrlg2HSbxFTMNB441znKrUFJ
EZ52TjxPeZj5IPuj/SwQEFYDXJt/gbmdwbSb5QccvFYcupq6iclPAZcKhNAVN+2gtS61MtObSLsS
/aLPX98TCo/u+LD6eusS1QHFD5QIg9bJjwulayxIzShr/HVkoWgriV5g8tHN63IwzSJSo8igGudy
TtEEnPKZ/x+k+5tl73n+yDFUawnBCGEkPjUbVHF6X6CxbA/tMbdkoY2z9l/UN1XNgulTQbmrddbo
jVrS/daQ+szypMzbIGdNSayinyjxnYdS1xhfJMJeh5rxtBgJk+W8W+gf+nDKlwQ6eH6LerFn83ux
oT+jCOsHKGQ29C3KjwoExzlmNqQ9lqVxHxY4B2lWC61AnLLEzCDGAGH1kPUNy5W6Y8NNq2CgMlO1
ltReXHrICATqK/RZpBvVgIjPLuGVQmRVjguvk3LyTR8ODmbCBlLLCJtW1Wa3sw7pwGNXKSm80f0b
mT/U0f5VnodbOXPXWI9YoAYRRHtIlzdCMbW6mW5cV3Au3r2Fr41CsE6TWJEmD9TXNSmcRswaZpWE
MDUoDutM7sji84Q48aQvHGJBVSDqYfiGVzrPTDpSd94J2aH6DnWUGgmR3ues+bEwAMVGs8f31g1z
9vt+RLAMf8XAPEPYT5xghwTID5xsQhq8VqM7lbVw9XK3DBCnU1nWIEmJdqxqJ1rvh5IpoPDk1HBm
D2T5TqvHaiU2NYMZlINCRynrXIjEw8MLVhz0yHNAadapxxUsmSM28/TUkjNQq2irNK1fcWKyplir
IxRQsJRLNc4iNwGkw/2BAGYBlVLrsMYnqMnqLCboDkpq1PCvQU4cAwgv2cnEkKCmz8a1S2Z3RrN3
cnitRAPJUpp4isN2kxg4IcSZQaQR65XtFvaPkXKliPrQW2MM1VRyKKCC+5WT4SHu5RyFD0Ka2j7I
8W4LcN1ABx87n9Xs+JrYWS+CkoV6x3hQWEL08HciZnEz+WNadRcyVksmbWPixTarm+CfqNZmgUyU
6BZ2JqLd9FHDpAwmTxjjiWv4L5wLNXX0nrAAc1x8pdcOHi6df8vorgjyj6Q0ItEvPJlsTSBhiW2q
z+k2yxaQQnGE966UIBmW2BCJsAKFxmCRaqGuvS6hkQjoerwTJfyFhuMLuUIZt97xjAr/l+GXeJGB
4iWeLnHXHry3ufRUjIGMdvMOK4Yqr/seUIl0N8zRQUby5VtJ82KixP9wp+85HKZ4uo+Nc0YKiJqP
Lz/1d6ViuUPSGkrp9/BpxAvCCNulVF334LAxit6++P+ZCrEycUY1K/iSPdNhBNX9LQKOlsO4Ouln
2Fxg5hXS2dMYQjA4IZWqdi3owTCU+laJ0A3g9EX3RkdTpzzY+fIayTUAgL71liaS+7ct7eJVCGO8
LF1T5dD3Db0YgVhKhLEXjE/VwQRGMxcBzgA/Q4x8fT61ndaH5oARxftDzN5WiRJgW4lCx5Ik7HwV
apj7AHhNUvAV/TCFt6wunTehtP7tQO1Vbkee0CYbUC7glpYLQhqP6uoZY0IHxZSzPDcrRzkfZjoT
3f0s509nsPUNHO/CVyNrI5fTxI9Jy9NlVQXp4TflP4VTP3MU/QxAgiTHvxNwlG/XoSUf0xpnMM/5
AdnhIQXAMG2bIgkNR9rjVzwrknh8kP8ajkYXKbSOWR32Vhk2jhoskn9+EwyxqHHHpTxVmFngrsV9
sg9nbdgekmpa1a+eO1bJ/n4fIsDLicsnN6GRYd26oITeMj3YWH1X4gkCnTaE0oiLlOCu3TViMMy/
pssI/Czp/dZldgUMKbZSmbOYXx4H1qulYzswb4u6diSaYbZ0HtjHhdxT1otOElZ8i2XE3B3tQ50e
oOlC+7nDjk+321p9/cxCYVBqpVc/wt1xPKAECPUqcy2QZfBAXWmtC6E/kAGxXemxXuM2W06KsjFz
LwUYoQiUBMxmXuFZVBbEDjJfzpXKAQWkyipQou5I5hhCKvFJUavI83FvF5kOD5FIs5k6tG9Rr5Ei
SqpgtEij4MthZJxNgUdjB9cIy9ld7DPN33gYE9VpIbVKx8vmTnWA9X/Nk5a2GlbJSBESTIlerbai
8o3ju07PQae1DkDbwlI7OYSfEBDRNFzuFjde0o5YxEjjovxq9w9BYXgqdV7ShnTbJzzhU/SK+1Hx
mTzTsT8bCHvqN7gyREoUg2TwDTCTzli2QLEPZuShVLYQHGdl1rMhPHcmFpQGmBL/6PxXIDCHv0Nm
xDnH9ovB2mkomUB1aguSLhghXie/PhDH958/CvJwCAsS7HUytaXhTvQIySqXD9XHJTcX9QEztzm/
8Cdg2XddZrz3V8kyH4IpzrP69N8FGBKL4A5ZXvFOH1nhQpiGzceBbIE0o4zehIBsQqOiiFpyIOYa
zwWq/dq21EY9X2YEjzLtu41shjZlaV8Wo8fovU3SMcDwiSkLJt6EVPDuGeHDEfZAQeJrXe/8m0pF
tA+KHsMyW4w6LQaGBixD1PPNhRh8F9NqALhLROJWGXXK/oS07irla8zDQ2Ky+9KAku5nDWVkfyPO
+BciYIPD8YS5tQWGdBZCxzoROkEF64UheRSePfhyyWs30ZzGAAoqG9H/nYYJ9dfGZ/5e67IJJnCj
oEK0P+oHddPaBv4+vGJ47RT1a7JZ0Bo+6d145hinOZCKbX3gJokFSYXZzvWmLsV4S8dMVCBhegEW
tybGc4YAXTS4AOj7GIEjfxk0+53/M2YFNh8QT54Cc5rDE118BSd/JwfPFA+etc4M1BgbauIJiC4B
9eMHqtoXCIdFVmIZe/Tc2MnRQticsKi3u6bDJMkm5QqYDKps8STCMma5oRTWz2O57UGDImx1uN1M
dOo3VdpCefM64DSYtWjzfbtrHTtWlJw8qxMlMAN+YxENDTE4+KXqW6JRsvAjlNrYubdJw0M80bLm
TEidMtt5/7Q1OkdkxDuMgj5syHxoRTGaEmSGzyzMOcu0TZP1tt0ydmcuS3025JPNY1VwufomNEkG
s/rtenhjzqU9UpDuSpEEo9hysQidSLCT+F8ziH262aLHz1Rq8k/aS/7USmp6slTxk4i3wswMThSE
mnMj3F+1vgiLgKv8uYc0ns+tJFBwj2nrNHUV3b9FO4cVlM5O4Qx35yCJAYMF7FtAGpqCR54Jyx5P
CQ6DjfhQb8PZy8QtgZG5YjbbC86PftoKE2Pz+fCer+IaKc2WpU5c8jeTx8iiQ7hYGznpJXcRwhyH
O68lq9rtDjN5qua8tGARnJTnkB+kxF9zZ/tqv0xT8p04JHZh16GjSFkXNGgYQAb/Et0GPo70euW+
XXVdDFienmKV3UNAEbnKnY3zU2wn3Z8Q+Iek+bH6AkpMN1V+vy5MhMcI73Y5fwK37BIMilNqwW4S
W2BkLHn8DVVCa+vOU0Y5rw52Jdh3LidI4CSlBqTiojhaCoNymhNJuoGKEfpkM47qf9NPhFBNeHJk
ftHV2qjKhf1EZ/wnzSa3jf+Ipn4TD376weDf7vs8ZWK/nxILXt6aRZRztdZFNM4CWfwSEcxr6t1R
p97Ze5d0XJEUMH7Ua+kyAn7kZGsi1OWjdtCsXXqZCzhldHpdPrtEJ0PKW4djdZDJj6uUNIEs/NvA
Ets58qHpF6HIWIBLVB5q4cyL633VnM3xZAhfFhD2kFi3apC+easI14llFf1pYJV44I4re/xzU8d/
l0vfNA3gkVm/WZ/023Igv+CutnbndjSceb14p/0AM0MVEu0BfpUuo5vKbuGhI4+UTAXG264Y8var
lN7M299xZP2a3uLf+CGR4GMUsM+TuvpmnnCjabB0C5hYqGb/ru57Q/iYbJZD/SnUii/DAQFS5K3p
k+MAKljrV9m9oy9+zxFBNYcYmlHKg4XyLZKsuhSI32Po3B7RayOR+ZT9Ie6YhayK0aMPEZ/6TjeW
wDUN28e9xoaRqamxRcWoNQfFHfOI3OzrjlW4wdjozQ9/oC3JeG5NpcuAeQfxhDxosviQYPGap7G7
bv3WNtIEf8E9rxWTUIb1uwgxxnUwvtOg+KnR6IlReS7GLrKwXHBP7YyzSOJH5W007Cjbo0rc12nd
+R7xEhT5zaF6gtW3EDSNdLxml3NTuKej+NcU8PIveCbCauU12c+C0BuEkg6wvufBUkArtrb3is4U
f+hrN1xztWXHjBQwdqa21umEdXhgkzuGNkL8fDSIxBC0chpejvrIuvawodWJDu+ZEGcwJObUjRAN
YtSu0oJVqKYT5OE0+myaA60x/c4VSKlK+8WWpFPSkaOsUZxV7f2Zm7cqWlq+FBk5LgHA4WK9QuJN
w/I0fBnQxg8JqbZaQWhCHv2tzlz1pY+m9jJ33yFEY0vZtZmpMwIl0XSzy6hfzykr7VwuysRCiWYx
PrBagNdCRkzRg5BKdDsnuG6C6DJ7/7pUC5GV/Ka/Rm5Jh0taspvP/Vrmv32C0nEq7ZYjAG2Pswns
8dZPBld05xxIRZxnDK6bcOxOvMDPSDG7TUrKy82SiAGVopkEu/oULm0bhp4cJ7gJPCJpz0CmvS/r
313hsd4d0RnM9NKcMhTOxt/odsd2c+QnYYx+62tt56v5x/Ed6K2XnBnLuBeAXCRd5oJmigQIeRz3
/G5KEzp/DXzzzB8jQoaKOibqSIEsPob+q9Yd753VBFT8TG97x5QIaxxSsysTf268RMiPfXTHywSN
IgfNUA3YlSaTEwRk2YcyGLBic1ZEtfxOCRm32ENAg41fhxB6BJc+U50BtyTnRAVa2VGiUmqLOL3d
2Cqx3zgiFlLcdc8HgFFqvFmAoiiz5MBf7feI6vCfQLDLko973GIZgStVcR7/jFTiOhLE/pY83I8k
WjfDCdXW4wqPVTQE1yCbik3qucXZWtiNWUlxL7+E8sg8uEV+mFcwdymLFeeEL6WK6IQv65PI8OAC
Z210E+cPjmJQ1jwq90Uf590AiZiPa+l23vFpVJu8dY0khY2YL2dhcXdktqYZd/SpLejsmhMLODBj
Ry9PHxeIdC8mchAMnUL/AAM4W0EHwGYx+ShvmkjvKXJLWQRIU+XVB/Cs4aeRdvYItF5AWX62icHF
0o5XUtYyBhv9zDv3IOAk0IROHZA4ClzZ10yrzWsge/XxbbMQnA65CjMF3XdVGrN8O2xXHzw3Im62
A+x+b/Z1C84epbkA0uMgeM/KRb0ZCOL1B0vb2EvrUlFK67lCcYe8UPFzJ7LER+JM/kcfAGz+zsDy
WIw1XYjCq7eDiE4EEahFhb1SFnTzcISLzvP99glk/q7zivKy/gYZQaCvmKEJH2OXEP7vDYg8cafp
+l7ckRxol9/X5vaKuEHwNlelRFeW8ZfMUmAqa9qvV1BQABbro0LGbBLfK5FDpbw0D0BMOpLof/MS
eeflXIgf2TOc/m4HREbpv3YaBjRJ/0JsmQ0DaHmYOe3OHmgXVqA041w2f4D1wyVgnE+cPxBIsVJC
Epk/o9Hyce4FsMunFZFTKmV9E3UM0kQ4R8QbQraK+KTWYyp+FqJhKu8wrDxfIWIyuDNp5yRlsSb4
X5hncmWWJPJGfnieXZOAa7XzfZvuONmAWLW08W8p9cDDL2OKkG4xhdUQX/KNlStpW43zRAjjJIYt
vjZVX5lmAW/Lr5ZM5uN8MvL6BpAX2lo3xZktZrmfInSv2qNM10jx74cSUJ8SoeL3oOaH7KpgzMOQ
pc0167zDj7jS5EWXgfRFiwrLrlnd7IZ/m09SjPVzQAXUa1U5DPQLQZYVY4qFv2ZizkFLtHlB9b6n
pjex0Gje/KbNVbx8Cr2QLlCYt8OL6NrwVVfZL3LaozVwVranIM49lwsSWqMLQjjBxJ9VZIZJ7oty
T3MYRz3Td9TDAM3N0qTiTaFj9JGTK87xvu1tEPN7fIn2hLwh9PbqOySAQAUIeWpzv6kr6WdSNUOq
BWVlaqmO2l5co7frp4NRi/1OOCchCzt8rpueXx4Ra2TsNEySuSNKuBLJ1XEWL7opOtikgQizFZEN
8a7Ffcv2W5oUGZuXGzUerDHJmB8CmjBRpAQW0fUbjnKyyYzpFVwE5WtZ/Ysuas/ylQd38oS4MvXC
r2y/k/K6reQwNuxtpy7e6JWKtsfMT4KrJCmuH8GGToWOZXChUA9E1jhlYQKoZNBrvr5f6OsH8/Oc
URCweOtxXooEKIcG95VWSftXV4SOYrUyaUKvfsiOL6sG6RSG5aK7+Q94vCj7XsYUEZV49mgOvxzT
kcEO1tHel9oOG9fFbedzBJWtdQypCsuHAIKnKR4hF0Vv2IqeXAfVhwql8qnb9lRwebGRjvoto1Wb
3lbgFc1c2oq4uAxOcIb3BUMc9/4Ri3gnBheGwYMh/4EDyKbFW7HOSqUzYf0MD3kLeiERW7TDc4ck
vCC6a6Maw+/wnyKHkMaNJLdkg3HJmAE2TQeQJ2bhWaYKmNky3MZQ0hgYu9ZzAIMCA1uLqv5oV7en
ztRAnWTk8fjnAnMZJH7eX5+StKFKHLIRzbnfLNmhXgWkutLq70YxlHvf//6LFd3oX0fP7AyFjV6g
Xvz3P5vFJsszJEhsYWifxepS6pbhMc1XnQSl3CdlUDbK1LT2dENvz/fn7lM6Bx4tKdHfCZZH5kSS
HAl2lzvExMnFObTNC1c0xTAKqRCpHbwdXyHu04ggOyAk/2Z8w00xbvLa5+yQwjdY31EVWS892Hzw
z78nTo1MYRVysTgLrscf+nXIBaX3SAvFVs0lwt3A9EhGO8GIywpz1weWp0IXqbazKS+iOM6wAHTO
+q/2QNo7gYfGnOAlsPFFuh64FnvWm5L/jydyI+PzFcfpj/sshEMniap0Cfu6ZVTjDFj97u9NeKdT
j1S99Ekn4m3rlWGrI/1YFV/bGMydEv9Kj7EJ0KUQq9phJF4TmPOiqY6+O2rUqRrY0ob4faNK/AYk
7ZzfxTBsnxbOeQuueRqygPi5eqAPgB2tLudV3QMyEW1t6DJKIoLWsih4/b9qQg9tttRxEFYJmKNd
RA4CrS+FN3PCWIiP5o7H6jI6iUASzsi3Fl/3AiDyq0YYLHZ2MYDk04XtAESnn/sEyWah1zcW/5cX
e5QqEw5F8CgKU8MAwcGXOmm3vnxcAdRclMq3rGZdpcYBCax4bXDFki6VVjAn1JHi3c89O5gvrHvK
nthhFEHGjUFPBUR2pTAgW/VvlEVEOXN7xFgNNTtmRky9loor32b2WzPQjo/zTQqyirgxubIAv5gj
YcXOyl1sJTHI0I148PMJspJuPX9NsT+9hKk5grCdkQ5hawHpsse8txwwy44qho5sqOV0dHcFV7B4
wU0mV5k1BgF2RcQfy8sxsX+1I1nRdWSnhxIGTVJbtx5FeIuOfnSzxoAwFwwWnt+lwX5mDvQLg2Zj
u58lv+8/8U41wgdn+y87ErE1yfRUfe9AN3fsAiemd1kyi81HFlxbGK7x6okls/9lLR1/gftwuSys
Q6N6xWElqApj/H+naImEu5evXukxzcm1i+6lcCv/k0WRTID6QOzYg3seS+H5n4xlxdTUv83fJxAV
fuhuhzn9RWyVFiCbaAcD+i9mXeL3r7UEv6xEn7DuXCAgh5+bp6qydbj3MoAvGnAgxVnYO89H3/5s
HA8SbZd8M3ZrYWqmpoXD1v/X/u2ycpzrw5fsYhPQkwyKojJHF8vt2yTjzH/FH0i2/m1J7CjcN8Wk
9xJKT7zMeg0VyczvL3RAL3JBdqRzJtej3mhHkAERAarWgjB2g+jk035a942+9MNFdPfzxFy7gLl0
/HKAZRV51DQSMa8u0d6aNGChxHr97d5uKml0GFoUSelpgn8VTyfzmPuhhSMhqgJ5osUTOxsz1ZPF
rg622idkJ33vmDmOWeLMxZL2CUZRFXWP2XzvMOlE+a9hQla9wYVX4sEI5vbZIqa9byx+O0eLsXIo
9WQuc4RmspPbtTm16phYJWvfPgAEzHckzTXXZK3Lh5bWcyXVDWPLAsiTN4Fsak+Q9rK6sBdFYhVc
DSqDK1iJPEIxjEIKGNXfXxI2CLEoMVeIQ1EYpDSOvL7+Gvw7yxTsSCUpg0mkD+lsyNJNo+/DwpIW
8Voj4HcfpeNG8daGDX+QwO8vfM5/ZGZhlN8mm/CJ3/Ik4w1punTTTVvXKnik4L7TBF1mjZkMEQ3O
OCAuoPhozynyPU3n+nBSCofMfgvvMp9H5aH/MdPYBw/70Cn7lDfQaaMIlQGJ3mKYabGr8vq3kdNA
liRRmPn6GA7BQZYwG/k7jAbAclaWxU1etfY8/NbOIQdvDsSo1qGnNzOh6EuyLC0l2D5iStTxp7wc
B5a9cbeZWx38yjZ8f6pCqtVWVuWMUkvwVoJ4y0l2FbWGseBCBaqJFJXWu9ylLj2zJ59sSY8cgdc4
QIALvCtCwM6qIKo70EAQcvXckddSt+YGzoYKl/fZa/yHnaSkrEwKtXa8zm1g1ywguqEwwLglWHTT
fedemPX/W5NILZSUxHzNDukwrPXzQZqElozcU/m8ybExODP7rEq7DjxLCPvbE3HlpAzqk5P+R4PI
wCrr/5aOPA3B+Fcm3Bw1KS5KFPUJ9DpARPkIMOH1eTasfB3hRXNJSWvrTEYe1mhLKzD5cbejwZAc
8wJriV4cSq4KatClVq4v5Gj+ZEYYm+X21jNn108EXNx86oNlD+5ULelu2t1a0MK8yoTAmSfH1BYA
1/CRX8ATZ3J6wTDu4rDPeSA3ZqVf11ehmRRLPH+qr+Eoukolh99fYku51cQsLAu5bL2OX+CY/cFW
Yr3wk+7I7AN42gT/CtQFRwb8j64GCHcNHxwEC/srjWWqpvdMbW/ryrdP2nHSfB1PrN9JX+u1i27v
krcPKkxORNjVNoh652vVUeM53JVRyI0SukGGTPueaMyQMqxxMR256jYlZ5GWwB87gILoMnT1W+gM
MjmverRAhbc0izljecmYPZFhxWYVH2QRYnT5jIqZBB2v49l7lkL5aCScZ9OFqH/1Dofwp6o/HwWw
jcmTF01b5LPVDtvIOaPrYzaprIDYzWbDdsuGCn1IxsPmRvEhh8C7+58/WTorkxdWRsh3A6JPxb6y
Hw4OiGJSxsdt7q96QaNda2nSM1PmfpK+YNF+5kqVnWDNsyYxfogd/hJEUeNgycL6oZA4reQhus5C
kiWkW70ZqE3/bhbSNvUbQCIFgLQNEHYkvCGC8czElG3KQqFUxfMjeEmTsox5J7dzqDOGpspW1Gir
nb8LRABDkvubpKjn3MnqZ7w1oE45FrMm7fQ4nQSdCvgSJj9KtqqA4o7SECKF/9ZtfX0m+nJjoP94
LjoCKo6P9WVxRO625WEGEkfHa+TnALXElgRk2hiU/hkXeztCL5NVaVC6vMjUXDqqTKCfg1O9451I
955NcIQUE7GnhCg/DduZB+V3vbIIIS6TBn+JCvzHN2UQysLz1AL3rSaNmQR/QuIMj7gXcMIdI6rg
CHy4f1KMp1OuMfL/RSh5p08NyjlsAszHmwMlWKWyzKtv0x+5YLWttolMTbZfxOOJdfHD5Wd94zIO
nL4N7fePtu1A7JyAGLK5WyYExyWip1oDEBVTAenuzTD623vLv2HdKuX4eGdPYq6tKa+mu/e2eenx
ZP6LTjfYCLuPl6CfAiKGkQww3yfhejs0V/rRq7WXOV93bRUNxWtvFR0anCRKVDiKSCOWEqk8bTr2
APWMSUaCNbytN29S+WCUy8j6juPDROGuA2mMnojwqANWICuqsYm6Mzf1DYG8RezZvg9adEHFa+xV
sNS8GFsImhd9vUHpcsBc3zD3ILZJzjBMKKGMHSN8yd/GZmRQ3mu1qIHGM5xr5zb3dN0vc7zJtg8S
GWnc68k8H3EfIfj0OllM6S+ooBzI8AB0CFmgrKeHJ8wDgQaw3LOI9dA7NTSVTuruZ8Y7bj1hhxxe
g7n7syieb7nzYw0aoqoq+t1bx75BNpsVekzjxgKHxtz4e0StNug7LA3pD/FW3aczyrNWQV+nq2cH
yiMw79T0qb+JWR+7Q21Nmh9Vmee0LVGO6PXbnX27QZeGhD1GQ8rIsEPgrC40bJUHxyfG869aD20H
qOEGI2A7f1065CjYolxzatmeebEeSqs6szXDySwMF4BWpg4xiRS5RA4eKJZoQp3jhSR2K4EbybF4
efCaV9507shHgKQdh5hUPklXgicON3ssA3w4Wu56cjz78w0u2pMVectClPsweQKvqzy0AWs1N9MA
3D0B4QkfiLpv1afcG4N395Mx+Q/3DL9L3j5aVWTgLIXMJXmofmRbgJR2BWmhKNQAnTnMUjJXLNlz
YVMLVqBxm3DbpM2UXqke7HIul8zJlr4V95XcjcpAL4FnQBAsGspev5i+DMAkxSLmoJlDHb7BcdbE
Kts3TCrTWUO121viDnUrRxUu82DPxDfkunUVu0Uzvzk73qogW+AriHwpVFiwhug2vl10P1vU4DBS
usi5BRTyxJ5RYnZUr1U+BKsiZBloZfovuJXolip4umIIsfi/xzXn8/SnLr8oNc0Uorn2nS4jUFSF
DemOs3wMPmDwrGJ7Q2JhzT0Q4OJ1ipqCuLXCS2F+k7jhiZfBF3FZNj2NqLE+xBmGFAd40hfEIvO+
Bk7pY1z4R+hxeYWm0PQC2BMcIWXbrc8bifRONCVyerLduZbKCvKUWxAtnspqnn1ki+WLBwNW1ZlH
z/+0ZxILtaGjeMrqZRTy2mqiLfWR9EUSBmLpUOdd54vdhTSCN3AidVDoIKMyB+UuoyriFAsxTlCl
GUd6l6xUhtN1djQSwdlhZNrdta7JqdTByNSD6AIz6x/hvrEonFK4DZwVWqAv+TsTDa3DaJL/sRJh
NWidzhDootbBnLVA4iz59cw1AHy95IbsFvLg+Vxk2OXxkrxTvBg0Vh6XWuyM3n+oO/FatVRzg1Kz
pnXHRU0F93luyBZ44wFneHdwHbX939SI5FHFbEDvaTDHw72QrOsQ4k+CQk2PQ4eE6M1Gd3yt8t/s
dgbBs+pq6vkG7/GXWXOHM1NTpvEAzNBdWGWuM5YG5qemWAvKnFK2CYty0G7uiA/KqbNstkWgLk5J
gr/7cF+ipn88DTA7meAjEx9TtfV/w+lfxAW9/Uf5xWBv9wknLoqdWntYRkZ4eJrz+Vie2Ju3WoHL
cFNiYLkS7AqdBF65oPYl8vWB8Re7AqtTHotgAy50bEe52MkHRSF3NXWEvQMh0SQGz3q5BoC8dxdI
soqZmv8AtI1Zd0k/JlqfzCM//jufkWCsAw4R9bXkVsn9b9GVDhxav/uoz8TEjNbUAzbpEw4uNYzD
v0VQQwdc2VMcDLucU6BJ2XMRorYPRo9t2LRrWwBDurmjLLnFx0GgjBsaRJA1M++ka1Jl8xPouHVQ
BR4sVG5gcrYJa5VRduZoLGx9QSaP1l08Y55odcDVS3kNPbHb7ACJvECbf1uKKocXUybyKLGPoOqB
89zKbfHHVcSJFjpu5UYWGelPQcVGxobbYcRN5d8ZInv9tjQH2lI9KVAjxPxNFvrYYToT8WisU2CD
zAPVrv27PtaIgaIWNev12m28xp019Q8tXLUzA4DLWI1GPpsqzA7ugDrI2moNgw7blfGlh9w/70JR
4g7GvM1KoaZLNdIjAxZhtZ/97pI1V6U6+5wy2eBRIJeEILAIseeqF12dQu8ODCsFxoIgq9ZGuEG/
79HjwnXOSVyGl97UgGLSj6zKNmTz02Ca15AUxCu0mgJhNZG1vWvKDQVy6/kA6fb1lktoaP5wWvd1
zfjG3b6W36oPv8PyaUMFyMn2wh/EwRGpeqribbhZBJRqsqszdCdVEd8vw6fu0JnKzMAOjBtYdcfl
pi/L0dUIQBDwUuSGDTRQu/E7MejKyZiEVDHj8CPVUFYV4WDdcCcTHDLvDfU3QZ0qvhFpKbfjuR4x
LVL+NPsyk59Uu+ae8yV4iSOIHNGxxYL6mq/MvWTtYPtNbucZz33iOfde+bTNq/7/ae6TX86KxImd
SX4b8IC5oZBah6xOJGAmubNRXvyR/ukBXCkEYTJUFoVjXhJ/4UFv9bdjFyMyAVKD2PnbU8U1YJ5s
A7YQhzNg/zIUZvd9BQLOsOQTAIXhVInDo7I0f90jC3OGETm+q0tJzSc45OLKwv5XkSq8GHK6QnM5
7GuU5Wof7rwDXWTWSNniOJJTg1cIIXaoQadp7LgyBsidArbVA0lfzsdi6aYgMZnURUoCfZaUEiFz
uLg0/LSsYaLl4r4QwXxQlFFksN0cG20JliI3/vThzkVviMK4PnG56p3Obnpg/AAmkWzs/bObc7d3
03FRM80JMRSJYkDftAN4fI8640iJObofII4DdP4W0yTPAwnm8ExqR2KwHFJFL8ZqC5xUxLw/DRfV
szsEmkblSKi0tMrZECCEBjJxx3GFK/RstAfL9MzxS1Ue4VM9peWvzAZwGRTXMeYSK2zHi4yjIGLm
ldt1K3ZnYWaDME5eAEWw3sg3HUyDxm1gXS1iS4BGzszb05IuMgW2BxcB70jKjNXZASe2G5ElOYar
qZ/6bKDqbh03GsPHH4lmUNQ4vVq+0N0kXJZLtRqu+H46oCfSUDsIbi/ugXXR87jBTfhMbT9XorFy
OLh9NS/S6Bvim9Ozklf4NvasC8BTwzP/L5hUF+dhi45Z+T3e1wdOzqk9VHLQhSyeiTVqu45ymFjX
YauhVRbFlaZ5GllLc3+J+sCfjhGqKotUOkltIJWA5FsG41UTpzub8JhRCzESwwDp28KgXokR1In9
16v5oeNpPpwkGsuBIKWclFeKKInT5RVzlGeY8pB2WvYKlh0uxFxO/xZ+oaZyz4VHV+NBQdJvjkbF
C9WQSYuK/21pA79gKiKc60sbojMwxQ5kRxV6XGHFJuo5+SBj9Z0b0+k8m3VnbS8BVlFLU8ED3ubQ
RFruOTW3Sb9JcEow3PgryGuyRQJvB31dWyIXWWn9CzqJEToDMMfLA1TDnsvKYPVK1pqCA/KOMDjk
sBUh+I6QPv/iEtQg6qvTz7CNWu8P5jH8f9ZgG5g+7nTfX9xGke19q6XybTiCp8TPlqauEVGSKJ0w
VctB51g34I76kdf506aSONiYuAq8S/0QzBu+lCXU9MqoS4RjsGP7oRCKNHWgw7B3Q2Dw9QQwrKds
U4YUxpba1jKAJkr4uBmff+U40TV0ODlQ1r8sJjBxwexVdGYiuwAtr1NAibT8EfL1pqJTqbfFZ5ZS
s4g2wC4zJzvYjNQx2g2qOHHjCqf1Sa1Tn5m1LJi24XI1e5Rcgb0r+ebAsnLf7p1ZVy1pR59xFbjo
bbeRQIDCbelIPHbwMAV48rBtI7f12m6w4MYE+k3EmmffDu4crwalkb3koxBj/ss+8tfMcngfSh4q
dRp1LaAXwJDIoI3tn8XDWIgNtiVjRE3vHWVmQBjm+UJ3uXPweKog6PD5xXwy950NzVx9+f590kDA
HzwsD0QzYCAdmMDthz+wZgfR00FbjttzI9v0ldF6BqwLtDTKLN0p52e6yAE3vV2vuf7hJIc2xSZA
5TCn/5XVrZ2Srhbe0/vXuK+NlgvFZUDyU5RqgSFdahTb4eUB2+avgZkiXfIjFJvxHxp35J5l+KYt
Fy2Es1GiBuldyCCh/HYQsyxAe1TcN+P/9khbjeAVcSCAyVG/2mgYd2urVjt/zHxAsSqWxLWSw88a
rDlOZahVLPG9yAdqWXHQjfBsUl3E630H+nzNHAW/oRoP1HF3+6odlbwgnj2s9bkqtwCwVxxHAlSn
1EjUjFCMO9wrtRZvm4kMNntInGJqYYgwkcG44fPS8c5g6sDHiV0lUkaVFLC9YNzfdTIuJ88lkvAw
F+/E8VQffSm0ohupFp+rWBfW1HlmUQm2sBxYiz4HOfaaq89a6DNn+fO2jdDyXMS/zadwhhIEBeKe
FIO0mMz6aSIlGTsijbKXD8mtE1SoaoJWjv8+aEvrfZpeJ8UN4JrkR2YFGn1ErPsCFFMXo2Cx/ceT
rHEPLqZyhtuHYYq0V1+GiJVWvEUkoIDv+KuRtRMiYg/qMVuEUrnSuAMnNBIgfqcY5JtqNre8x6ej
3EIhEolEkCGIDNs0XP9V3lKwDlp6BUMOkqJ5m1jowR1U3fHI1f5mgQ32pmjfZYfo6zVedJBBSaN/
0aughoGfbhMRrQ6HDw/QbwdIixXeOPsmprpl0Vne5YGH8Quoe7ANY1qwFqT9FBJSVvPc3u9WUCQ3
cmf2UKZBLv6heE3TQxIgyAnatCphCL+SSLsIyKKbnorpg9jjC037fPuVplg3o3o95wZUkv6V2lqo
KgzJdoD3UmcQqJm+9iFLiepxIzblm0mK54rhhgIiZaUTdTsPolwRnbMNaSb3ngKbCkoQZgEvY1Ld
elLUzwVffpJf/6UNmC9USwBXcpyVxLn825gwJckGEPSV6vaxS1yzgUkuH5nYYF9zzcehnF8P0sq0
Qv+Y0xdEGq/uRMc0b00JQDWbyH0DH/RLNVj3QL/3beXNaqiqOI/I+bXUWEGTzHuPwE/KZPo2Uz8B
BnFQJEYnESUf/gZrZRHV8+6ozysrKJ3Wd/i62y/EwWePlPZahUlDZFR1snLPQwXtQG3XkTFgSfVt
dLjsLpLxb5QLX6OQnC6oZ5NWeoZvrAoVDIzQyv4654JAqgHs1J7uyOn0FYwGK5r6qbx4vK9SHOrm
M3dXZOCr2lomvNtwfP3lbE1x3yH6i32bO3Do8nsmhF+2TjPHZ02sY8zw6XuF/yHv3sdCwKosEkDK
u3C/nonEdB/TwOyZxsqLouDZowKKJrtwIX5yRG/fkX5JmNyRRDf5XoIY0eIedWHxfndrpzYPwUo5
8r0CDXNFEWBxyyy5FoAv6CY3Z3P5+TbE2lTFwwIDEj9/V8aUZGE7MrnUc1eYalAs5+rAqYYu2ODT
XTmDcfyC+MIdRrI6TL/rJ/c4LmdGIqi5BTX2+zjiOfRRmYHAB/hgSPlSY6Wo1z+8IgSjw1oYgxiC
pa2ARgsxr1Q/S8bP0Ohvw5WLuj2+NGKyIc/nR+wBkVTewDeg+Mi87DRlkcP8y2QpiyID5oQzATkx
8dEMZszDwmayTDFxFpcsEdvPRoesvbY4pteN5rjy6+NeLpwtRvMbx0JLA3BaFttdr9SkS+ovJlKn
6dv6G3ojIAvwRzSRhFo+UFYrfdChiV3EYp1ppl4Qh7OeoUcECpqZobczOe98urRMIV5O3Q0MyEfc
EtKV4UgcJ3eKzdCyEIrdIxBGnlwpox+RW6FqULGzCY7xbNP6hi3NdEuIIhSudiWXr0RfLe0wovoI
xvsVOZLB117pmG4/dvtZoDVJc8GJDxUVAsr5VRPQdtVXqxSoeuB/td/kaj6/VXuctQwlZk3py2pF
HjFYHcMWDLNRjYY1k1C8B9gTbRsm9ia5RlOBCmqAVOi+VdpdKxVOXzQOH8Q7eAU/wWr/rsckebBT
Sbts7MlU/y7ZFvgsNuc9MwooXmlrUADSaeLS9JsUVWl+Uw/EWGM9xcmPciKIf0RNuZbFwCpJphZX
m6X+ETa8yoqirrB9gvhvzhA2Kqpo7y090YDGgfhl9vqSxGV/g6NTLi9ruOAcwawWyr3l0vJEiZlE
cMljJ2lHF1RRNyjBAZ/C0aoJwqWHWX5WKnKaAgt/yWacqwMof7OhOdVc2RpUeo6bJr2f0HNFuFHn
g5m8qWwaQ1Vx/xM4fsWRAtbuhWsGSEMiCGSAE+rE3bGGT1yNoQ4FZNh3hyo/eDOfB7dsRzdKClMu
0fbdgniFhPPI5xqY2a2O41KOdpxKvPW6AmV70xhQ7YFd7GIjnEKESmGEiLrz4JWgGF8u+jFKhf3G
t3TdK02KFjJjY7I+nSdATnhU783KjpyODHwI2EN6khbCnMjD9SQ7B0PmIvc3Moxvsywj2FcfAEQd
B//TW4rufqR3KObYon6vqvChImG6mVOCh3BPLFCCHERGUiTN+4/LDFJD9BPAwpIdv2a3z+6ggaea
OA3omTtqiZWUm3NJZqoYbyKWkXlR3HUgMAKq75lyLWYUXXNqNQu1DU/TfKG8QIqBqfnLpIi0aEJ1
WWVJfTPp78N0BjMHC607lwLgXM2aq8SYrBMy+OZlF4cb20cw/zpW3zmbwKFfQXLmk1kNNFqGIPiN
nRxY4nLLFrI2O41UCmHnuORavfAp2eM0M+ZD8JxLEggsiPisYXxynz6LySb6OGpjrve3+BJxQCXI
qX9Hqgvfmf3ned8PcS08Ri7Mvhwdseod8DplsuQl3Z6ujLTGQFFp6qsV+puH5a2K5H7zUdSGTEhJ
ShX5IC9alv4rxfMDupsyaAJJjTMXUh5U4sCpmZObUzfta7L8WKfhBuytoXy9YwbMpQ3P9SxmBKDo
XzhsXQFGW2sXzu5p6SMkDVf6kqY0yoZBThSywRnI5lV/FMuye7Bj+4uhytKDFWjO7T9QlutRp64H
15n/6Dvxfdv5eiFp1v7NBYWxLUa6TdMIEgYDgBcSvGmwd8Dpr8vH52Z63D7gAquqdHaxcPUz0eyw
d28FgbH3X/DiOzau/BgxxjnKHLlf1Cws2Dic/JV2an7HMevh0jwXBdW/Kbert0LozB9qFv4tdTt5
3tL6j7KJX30Nb8mgXGM4KbiSKluLFoKaM5Z9aFQleFNLO6nGdH0Jf2KJB2A1f4ccZll1NdEmZsKS
o5mXWEjDWPVXJmjbg8q+r4en7yjnsUvTqzCxTL9D+YyZe7Pqh9SGtbfm5q/k7DUeSORU/r61veGr
S6+DJ8WIJ9zuYl75EmNoS4FweYvdvcc8GCXe7YQIe2JO7uBCsRIPgN7O0NG/eqXwmF+p8nnbU0XD
jZq0+t67p9AqmQLfdlvqdItIFygSLpytRTfMsq2GAZpzlJv3DnbFoIshV2dhDr870gt1AFQUFcC+
tNCWedtVWO25JRsbt0EkuEf4vmqjJtt8zcbi0BeLUDYOlNRsO2IPgrSk02aabuOpJ/aV1mEGWh16
mpjX6Pmj1NoezKaCCaRa2WPIWOsoKWnoDj0zFkM7Q94cwSFvAEGz2FhtDtw1i2ddpNrbo5GtM0xb
Neefu/aYo6+YVBlflxks2mv0tu3sfBkGkWN+5mVSQo0yulkIzWtILuk2gDIobkBKjRogs8z6qOCa
xSuN1nC5o7SxXa9YidblJ1K52u6a70CR4dC/1SrIBPJZPRHTyXhxjEbrwmThUFv8ip+eRVPMr3N4
pk6T24dqQtz0Rg2i/gjaKUu5dCnN12hnHLmZijzjfBXz8+Hv4SyuY5v56xSytcvHIV6gGp57k71S
dMtSBLI5m//GlUhuMeeq7LXtv4JDtoqquv4j3IsEZOq6QfkNcZfP3UzuEwJC1dlNi7m2pxOJbII2
PH1es1HPhnwPefv6A6sy0ixi24nQOfcWHr48Eyr6Ey29RnjA26AD1AHQdOzWA3FWW+UjY9iNc14L
n0IcDA+3MNAXlAeF1YcWA+cg7jMWXW9t2npLwm1q1rmRf55NceGA6SVKAI9SjuDcCQommT1TY2mC
5JZoeXubb2Vh3v4AXLV0mr1NPV7qEcMyrGiRzks/qEeI600EztSxeis5bX1ZeIhZjQegRDlfT2YU
M3lmrPJbZN4IYqdfHB+EgSTxlbOJ9clchaHt5BPW4uMvOXPZuVpeusOZu3IcxXKSaWLmlFjWmlye
ixmJWntyapob8vreGPaJRQGsZbAMwiJC+PCQCttRie8a6S5UBmdFYaomwR2s45Q/BN/EMog7OfJ6
dJiC7sXXr6TNdGfjMXo/qXOk7VozmZ2RdfoO9roPuPBvfGcNI3x7Xc62y3NhlkPacVU8Rvh8/Nf+
OB6ullM4AbmN0iZ6hbUfYIgCSzbM9/UCwUpyux5+hU+WseYI+BwejFCsDrX5UXph2SeyfcTTlAQd
Qgc87LS8h1+d7SbKXMqMVyYtwaKa3gRqS6R2VHhAHLz+a7Hw+b2PrMknC1Eh6odPfb0lxmQivKjp
OtlxlfkHtlEaOslTB9G8/dRu3r97f+BL2OB8hF+EnxT0qQLAvPZ51P7DFCQuWOfRkkuXXp+fb4fB
/PoYJPWlNAHRsIe7B5Y4CzHl4nRQSIxf7uiHbialrBSCHE0uNjU+ZLAoGEpkD1+3SmBvTELN5vk9
20U1pU+r3rdlb9NaAtmk9wYqwYcph3FYvRVfzEYe0UDq5V7agsy5ojW0gE9kDs40AQCStW7w0HKg
UUdhC1ZggpTS7LDvQ1s6x3G0vBTD9/OQbRuYMCiq/HGCtIHJ+QPjR71GkF3UstLTYIIfy0LSU0z0
Li4UelriuEvilfpqj2G187hbRavY6II/92N5eZyl2YctSVXp/B2eKY9sSKkheOlSPPjQdSKoMHe6
k6HVPFrBpm8sczu3JG2u+KfwNdLER5l2soIOx/jKCZbOOE8b/5i/Obra9zjLGEQ0w6ER20aw5ulK
f02QPOYNWybfVwudbctQSHeJRURn8DnOcbtnMfcIpn1g1CNFxmztpSYBseLOyHyz6eBs0lWFZrCQ
/jkUrVrqyoqUAhjyFhn2e7Fm1tMI1esQAgoldR0FlTST/V6nP6nUYyz4TaG0ZEt0njjwYgGRikWu
RcHCnFRlTMQrXIvP/FMjHHOlr9h3t6RpUof/zqMPbB4uVgGB36k9S8MLhga6j/pTZrqTgETDui/Z
uXBjoOZ6qgkdlM9VzRfzmsEuto7l+sNyxcloE2aUryV4ous1cIfWbK/oZeGNGyMxg15bM/hI756z
P5h+uYKEPGP4Ez3ChAv+JWVW/8g3Ff+CiErVFwS3YspoPgQu8iGyvxUMtOXoTxoBHsNJjGAP41ZQ
1eFYEts7dmCTrW8GzvTAyqVONrxV637mHNDM6D8v6W974+kOWiKkE6f9472J8SwVcRMWIxf2ni8U
9LD5PN0uhMFkRg4JsgJ+oPL5ahFZtdkS5U7BHKkbLbYVnfeEnuD7ZNjUtctqkM9mvrR2KmDSE7tq
vZU1GyRlBmD5FuTCtnKAqyQxF6ON4a8rjUNA6AnvD5/159leTNLI38Ue8DB0zZ6FBFPOE2KxYP5d
5Y0sJaJ1Z0NAsfRpacivi2bZZaqAhsazsiDnz9oyIPMs124Qd9iDsrpXbXxMobE06lwN8doP1QG2
lxPLaee1tUOSdaIjg70iOUrT1tsdvBM5thvdPQYH98hVKpCcsCeq/IHJReCPfA7zDUctq0mI0f+C
vUQRkWzn6PIph/PWHPjL6IdYvzZ9Q7R90CI5DNjq7BXJIT/j/6Vq4bsXKYO1mYvzSkHjdo8dDWLP
b77smv4EuIv4lAeSw3A6Bi7NTAW0nRwHWHmP/3unzHelnCe3BIK2KTuRUliao2ZMwxfXge8CYlSJ
XhIrBJuAB2BgdgtSDZu8yOKll+JPL6iycZP73alPRj66QEKhAbZ+MwSnfS9kV98RkyUQLdYy0nvS
9yPkEwxuN+lCHnY4WPh/0IIG2I40cLtQFroLJuYSSjgb9X0+H9NuwzRcJb86vZUA8UteVZNFP7+i
GisnDkiivSedzOtS2pO8uimcJncwFeSv3K/y8u/E02Nd+WSSfHSKAy/sN+YTrYHTBMiVQgat5Ya9
oOq/YvOjgQHA0H9i9cxA5uY90qP6LUOXv8BSkDO2lMP9NfEwSoom7bLbH+S7OVbi+NTcTjnC+x6P
MpQ+beg/kfww3azYaOPDorUA9Y/Z20YLP4b693HXpOvZhdEdZY9B95tjUQKbLR2yt+gYGTCZJWOW
GMJJHxpSfydTRp8nXrSbz8HzlQQ/FU1LpTnjaufYS8iq080Y2NW+J66R5wvs0RyHWcjd/EYyfweN
uPV0ysj525DewfMswzUSvFImmwrlJAxwsAZ9eT4KO96CRkDm2rvFkNXsbadxyY2IGiAmPQyJWIVL
i+wk++ityJRMdM0v0BKBZsfH6cCapi30FC4cXKDDpHSBF/VrjsH/6YrHf0MBmPmYlEvCrkkMSAlX
uKDk3Aqex+D83K9Hc0OmeUk8PW1raAZo/fhXouGfVclB4lSfJbVQXwOZWy0emihtE3uUGYPCZ2P3
N6d8HHeIQgt6/uePVJmeGt1Ddt6aDVBNucdfnQWfWWijkhlcE2mqzwWUxxPbu8LE2geHJwQuBlWf
nrvt0hAeLppqXOd/KuunQtFfOpyEUfmMak2iH2rBpTzTWajikCya/VgxoeAH4nwP37Q5P50gTjVp
DSc2n1nPSsg0kM5E+0GgrJsGz2eGaP/A6Rx/vTuEYlWrkpoH/43w53UQYF4d37ILs6hePhuTGUWW
NUgP2/W0HbFcpbnCRL7JVWZeo2giDZv8PZJxbt93UJ/cfoMwGVEcmR1+0cstscKPj2Y4GBvzgjl1
smtags/vGD13GaCL0Cf69rH3msJfGP79TAAYE0ibNJvwtwLq7AyHpWl/fPu0H5+Buet/X2+wrHoJ
CvD7d2MqlDl5tFxezy+iWA7IvkktESLZPsm6DXQO776ebUU9JdIsQt4N2xGf7p9ck/JMYxnRyNr1
xgDYZjH9RfWC4WIVQZvVOP9+lEWNmX9vxegzRRT/s40Amf/OUjonEx8k/6AMsKJPN7BNCZOLZZAH
YCg1ddh2sLr5b2oiuxwJcQDwjspAgmFnzIrjnr/6gA9qcGDsIqU9jTERnYDkQtmYvMdDLu7Mm3yk
4ehvFQyi/+dnYJiYDWxaeU4De+nQ+d81tTrHCNy26GgrmWEZ+B5JStwBEaV+P9q02mw/gMeEOr1r
+JkBPsGNs086zyGpvB7/RzhULQn5aoQxaDVtg0a8iuhJkns/wAewvYJLhtz06mYDvH+XunFCy+k9
aXx/lHsjm4BJuSyCgv6PF2mwq2Sp/0fbTyLl2d7HZC6gVMALiMBQq3++oIsHi9Y0uhEHSZaZZvYG
EXlHVBmEDvhwnm6lGvNh8OpAYo9+g+L6Yr2ek2eZupqQcGF6AsyH2+sogRZ9OLE87WqpxzLja06K
0UBoCQjkTPB1fNUs9oJYg+oAaRbBX15V+LpSqJCY8tkVbVjiM4dUsctGC5EknZblzxMfFGluAjD1
+T2hODd6o7Qq2a7adeglK1eoYjReaRrdWJQBvsORd3xtEAHS6xY4elbuLQfqpINvC+T1Gc53I2/z
MC/T5HxLRn11KsUi3sg91xP2knCdLYg+vOpyhdsQnl0R5SOBYbj3xaKcREjdB+wqQ3/dcwuv3QcL
zYKKnTw9ipNKJO1Gn3c2M2fN/0nfbLCnFqTF4kyPQ6lDUJTbuzQXgz8oyqy+eHJgjBKcTsPDxPc4
HAYGYe9UOyQk+FaFwmfrYZZRTVSHYV6FQJkGze+jOS0qwsSwyCTrLXvnUmod4gjmYWJjE6Fl6awJ
MmpBpMLVAwYV9vuaebQrIXMxjtgsUdH9Og9z3lkKH5QIqRFj/fEYOMo76Bvjtg/P9obB6Ok2pfAH
rngp0MSDi70Y72pPaW2k1ZgkceoJdqjFHfNs9FP1Ealk8WpFtCjETtVb2WaPobuuVFkB9RsNJhTv
3wz54PAPvSEFn62gFGkYF7VjYwiCa8zAr24n4UqLE6A0Ssz24Nb3Iq2F5P4L2N2lI2L11K6kE8Bc
lhB/HtXv19yb5fokVXZEZovtKP2jmDmzvOEvFioQ4O2NanyFbL7C282aqQd/SmL3PFXs7xQnBplW
eHl1vBz8/fXLYoSoNxxxl/ICTk6C9tZVt4cb4Ch1ceFYAwA9x83iHGLPk+NdpzmnuSTnYKtgaRjP
SoC/f8un1Ya3UtjtFfmC8GXMKVuGr/zHZi8q9jGztMaeQV9ZF8B8Gfw6eNTtq7dqM8/Xv449Dzj7
gT5qb9RxKTAJdp0MzEIhXXGRv/zyETZHjErf+tkbzCtQqQ/P9/yNiOUH6zO0f1u9Xj5FUk+BuH6K
xk/0qvIUOpepRCoX5v5ri+FLbraPaMUADhmL6Xw6OgdKM+wEeiqJ63CA6BpzkPk5FcdAKuHnow6g
mqL2bG+NoyFmki63fWiQdnp2x7VlB8n1kN70qREJnAflL5TilFz9T8PKlLZJk8iJ5/9XIy8yEmT0
CXKbz6HrE7dcrHJcHP80LBqcv0AgRxXKzSjiAF3PqoaTbfcU4YyVofJ+FZSdB04KUmeRWnIJdSsh
szhgvONLUXhr3TWoqMrxpUzZjwXN9WOUh4UGIujmghoKh7iJs3/GpJLIXsPY5gSeCrIuAz8RAtmD
oKm8SSeXBvU2W9TQrsVnZs1HOFaSTdqRzcQBgorJpyajb96oHyg0lc5+sF++8i5TF3+lnCrg83Gs
mO8cUDKM2zsyD1Xf7wjiGyQm7b6G4sKEM8gm5xokzzBXelrfw8IbxdFZb3G6YgN5xN9bti4Me/ZN
73AjGS4GKq8XwN+cyUSIgA3c38UiAHezZqVuqnivLEjeIchq8/NLVpmbrPuKfaLnsLJIPmpwFD1a
MfsMtQrleN9CWWCyhpLv0c69iJaBbD8f9kpd4jSfyh+E5CqOJpAkfLSaJSSTRHcYGisn4AkngxWe
VqWFE+qRRMGW/Wj7PbAZAgfODZ4yi1EqHBDDGN/UuZAjyxVibdwSUP6LCfung/gpXq7+siwMjLIk
rT7slso6vBDZOM04mGKPJiUy2YUyhqbLnTyd635gTtn1YCa2pkNhpF1S0JB1BHbzcQpDQo+pS/TY
abN9sm+qCUNIRVr7SpzW6rqwdhbHiJqfcXLDPDFdU7KsRW+vjBHg4EFCu3knL8E5y2f9vDOuXUbr
ratoW9wrB+B8Saf6WtyDJpTeQ5iVePGhlW0j3kcgDMmvxHSWdSx5ywBAxDS3fWrXS5U5NNQ60a00
KWkRZ+oDx93rPWxNY9GeZKlAft9DyzhqjpPadxZ1a48dpR0/A1gl4gEum3/ZEIrgQ+x+EDMBMBS3
N3axhyThekOxqsPpQOXwb7P5BzNzDU6v5/klsCy2c2KG2G1Hk/mnA7CjDJ5NHeG7nAqnrtvKaX39
ALiAmthZEQMRF4RQGYVBkPfYkFvc3dXxydPQ+r2mQTpJws423KdxVJIf88ydnLxAbpanzttiU2Zs
lTiCkVJLABf9rjSURmjjGTVzyr2ysbxTExGvJGB0rxqmIx1Xxvbsf3b2+bF6+ffNfMaaDLVs1h1P
hgED86V3w17800WhKR2B/0uFj0JGcl7l3J+UxU+bu3GkfqIxZwIYwKG5OhrcW8IJRwnTKli54Llq
BWNQkxsXJnQrUiB1EyYf2+sd5uMU8BC7j3aLZWhzkQQI7SbvvYaxEw+GayC57aXkyRZ6QVTMnXQG
RAeG/njvKrNra9LVMfZXeXsw2Iml+n1XABI8NAqA04OUYgO+3XxuiytOew7ZUNX4EMvNe9UlQUY0
H63NrlzOiaCBnkwK+ISwwUQWtXF4el111ul3uJysRm9uZqRAnTskMRcZsIQkwzHKHixctPHuGB0t
QwP0zoOtPebpXR6qXBb0Fs9T4ELW1Macp8miCgZpHrhZZgmzdue+Wv6BK9LUVouTxfEJcryVf0CA
9REPSn3fzR24Lb5DQpZ3flZSLOf5ZUwurqiVRCfOZ8Thhr212CQ5nII5evfdB9EF88XMFAaIwXvB
DaI+PQXcuCMK3FAFgFjXSQB2hjkYKYoP+cqhWprCklFLforQqTCfU0A03PnK6d77wCdvL70rwLuw
LPEGaO/OoeCaD+JmwwPwiAXrw2+QSc7VVL2WZYKUWU9bMWDNd8gOpZ0dGPHcDzfRt3B8n2BzG4JI
HxYQfXa49CjpsWQI24N6x4TiesZPNKv1NQmBRF7PG+R0k1f69MTN/6KMQmqmNtcEEG5BbEUMDptw
VmfRBsQi5A0cGbpovF6/CCQTBF7qImMgQME6MG+gUZESl8x9WdAAvmmEd+We08XTN2c7J82uv8Gu
JCFAfTiUpSvQ0aHaGJPkJHHTb2y2j2k3nGkwCG9coxgiF9f3J2/4+qi3oVf6XKymIGhEnIRdSCtF
x749p+Ae1eeMHZQUt0H+rUE7k9JULC8q6/Tml0/SKv37sDHcY5/iQddd1Z6phoByu0cTFDP7PEH9
JBbZ6P1cWXvLkwyuQtuSkw+xjB7CS7dbVzD2CsroC+zG3VJ5F7t9b0oHAsocmBX5eVD73MWnQfr5
ZufIyzFfEdRt8PQaYTTUEFlUI9nt/IJri8cdKqS2Rxo/ft4lJZm/PCmTiV8kzHtarUhrrlv6LUNf
CKHZm1ZRAtlYQjxLAtirjT2ycXDwlapUZrYqvQHxssETV6HY40e9W6krrZoNS9zFlHoCR/Ur4XZB
kBI4gi5EwOlfehniYo2fFq2Z9o1SaKUhwreImKB9saZV+HDGmX+dq6EvY0ApNQ4GOFQqQKRQ2A6A
cSxBIVaTksxrvFu4cZOtUc5N0e1ezwrE1JZYjgIhdbLDV0kezjw4h5zXt/2fmxFRaiyhmpNyAS3s
PEc26zbz9qfH70M/OUZd6AiR54Dyl3ZoLBTF/dCU3Fh8HKBHlL4llTAsfh4iR1LoqAjXpVARUmQq
gfwLQVlzXlk85yI3MGKrjgmESJp29IvnC77Z64ffhE3Wvh5zqCDDOAXH2vDXXfrKkYoGELGFOXuM
2Zmvub/MOHDu2f4MWllyOqa7+GWJ2uDRc6j5h7Fa5/MSorAgEufmL6sLk7fHty6We+aR4lsqHtLO
wPHG5HKCKJXTSnnlw3WvYM1xC/x4xP5PPpRnAnEuG0W46SAi2i020TNcBiGZ9KH08bSFFwlgQV95
qMeVsQImvK3i71Tt0ErOKe4Ogbi3iJK1gpY2+2c+eVgdK1MMxeiJjRWupT8H6VkjU7fcJHYI3ttP
wUyj2YHHrcdtMAIrt+sAdssquAqGjjV2dcdr1vx4tVo7nfpwH4HYKkrEL7lMueOXORfydbEU+geD
lOrjYgQ8Z3twxu42zfCnBfC1koPwiScFPVHZqWjn/KC1s9mInMvd0hCT+Toz5R7fd4np9Hzwn1jB
dGAozAjDaz+S2ACs2CfhK1dwrP3+APd5O1q42yrmMDms/XN46soUjcmEF1Ss68REfm2AhtxvyIXg
KpFIE+oiIyq6eiwfFEdqlutkccNeDNqEASSnSpAu4GwlFcIp6NdtC1NiSPk8cqcq2NqLIAP9TWMY
CyrnkReRwHw8Sa1p9i//CSOs6Bh4M6C5DJLl8Vu7UzV9321IZ7jdL8+fM0qMPBnat8IgDBCutVCe
TMGV5k+qTl63wsmyLr84ism/QHPr0GeB/J0qEPUgnG7KHFo7icQgBTZU6lBCGeTEMlbVRo+VB7PZ
IMUbrUt5u6VPG/lj662J38Mz4/cQjbiMPGJdWgIVG1v+JTn8BVQcaoh7j4Dv0KSeVPBnJRdDHFTQ
0eGXVrOISXgE15gQYeUveg9/v1HrytbendWU5LshcN4mf7FpB5zm8LY/MJPMBFYGJcnZ0A7AeIBj
viFWO3pPzSGqK/ML5VwP0aBiEA3z2t4nkKYRK4TxSeFnw42eiWgwGE7AzPXWTa1jfNF5fOioANtS
JU3PVM4w1dwogkQ/xm3nqS5flbfOl0RQYjZYexRy2c2BCth47BHfgSXklKWslYyq4p8AbVKG8FQw
GoRoeIrGHGhf6nhwb0aEGIU8ddKyVp46OERnthzZK5Ps0DwdzbaBxXo2eqV72C1FDBoIvD7fPlvy
5pbSmk0Gsztoa2uYPZ3Qgjbq/75ySx3S6SijDHbrxpQZbC5RRbHcJqvDJRGHAQhf71QcmlMLA3QU
mt+G7ndHnY4YbOcBF5F3j2la/rtCQSletA/hhv2475CqQlGekEZ31tarPMBkoqyP5ICnRoQutH3V
AVV4gFRJRdpz03WeAwoJAdYe/3c2Aw9i8Zgx3iBYhvTys4XNFWoZ5ozxRYWZo42jRen8MfWZD9r9
GDWUwoWhRCXnBHVMiwHH03PvgbUtaCAiaWziUTDXWaEotHkNLWwgRsoWQUkpKevq/xCpeioeWaQI
s6ww2ujuGNjMyd4CSGjPtrbQ2E5AOZsqWcnCOF3QZSRyEw4iyK5nW1TeB/NO62wMpEXnik50AfiT
r8kDJqhIFwd6tAtJepS8NsiAiURSLjXL2dLUq6p/BhJGOolSmjG89fm/kDytwZfqGldFLHHo3+Vw
XPMdQs91iQYcV2TNDVsT83uENh8a1/BLJhZSHP15KEi4C1DGJ8XRCK6s4brVd9M4qXxfnaQNm0BJ
uS+mlySEj0IjSWK3H9S/LX+yvzAvQRaoctLWV31UMx/1ZqNmzY0NltfNoEXJoPDnVGPoLGCQQTT3
6yTxuUgQ5vzOlwEEuqrtyqJyLzOKppYTzaNNoubQVqoqCcuOMyALQ9RE8K5mTIn3NZQ6+ntVl0J4
oxWTeBIdKwvULMHEda30OVWyc+BpV4qMrEbLuM8jJWDA0/JhLK0KG8fFLHJ0nruaQYhfrGOy3e8L
1OmFnLZbTgmWBlZFhxSdZjbDzMHQL6DgiBln1yrDnYDWxYxZszyw5hvF8kwpamrqxSWHZM2sddvo
aazCGQO1gTFal9eOWlWT4xBJOtjo//xirDsgv6FzEzP1oMLQFfM8IBpOlSXhF+XNjRWm2Hoy+V/n
wYshyuh59REWRAzncYDASgqVY3A/oGoD6lQr9Q4+/nwqn26sN6uCza1oQnhMgH1kMgo7cUX5lPlV
mqun89OjV6oWBRzBPRRjBdZlxxrsJBBEJzLABk1H2JNM4nFSagUAy9wEQzi7AfOXc5ZixftseVy4
9wbhVuzdmU5uhIauv76L697nbhDwxnRwgvpL65ZCgXlbxfW9/pNyZgb1yx63slXMZ5Oqd1ASCyFL
9c0thS35vtAalRUFDfie0o3BLA2bl7pG/63wQlSFb11Ug1h2ratj+lFV7z4qbnFMHZn2ocQMyNRu
G9fzV2/njbkqU54gU+BYbAsAPQgIjw90hYI8nOHxbXSMKeyhPggXtW1dcTT3TtQTwBQ6bkkKRfAE
7VidnbQ+ej99c/zG0QVCfWTBSOcNHw3thsyUot/xRwu9irRgwTrFXFnGnejFXOutc3/zONBBibYE
e8NhLtq8+Cq27TvFAfetQE5cqhtru//R+37GCRXBBT4v9e5VuiIGi2Vd32Yll27JPyNb2o/Z4hDz
qZMyTW8/U7Umt3WES4JDNEwgRCRPQfeGQa+Z1SR4L9FPblvFqZQJiW/WOcS9OTyKpvJjbaux9U7Y
GfJTi29unwC2dTGskwguyODxq2Jdtne2Jzz+tD7pHsuMptcXoaf9jqPfgg8kkgaZv2zIZU0anFB9
NTHc3+gFmn/C9rzxq5ZyVGXNyiU/P8G0wxvHp0JnTNMXhcTyf5uUJ1fSE9KqN0/PpVuO9MJZ/qRA
iGShFn0StIDwFjJ2tzhC0iskyH8izObA5YKSPQ+jkqhywohrGEJy8K5ngfDYTsejDJPax7ES+9+F
pxqr6TlsFdqPPwx0Zmftqz26wRnpGW2eO3bYsG9ie4PjNUM6rG9574DLKqg5hZdeTKnr60RSHr5v
x8ye7Zr9zfWvH29pVt5WkNKpV5RhtjQL7Kk+G00sv5r+lrHwHQws3ymh5TyqqkoEEamNtE4HbLL6
wpKVdBUq44/BKgrkhiYpQ4rzPMwvEH9NLWFO+MDEPpDVJ1EqF+1fI9HETqYj/Pv6x5/kQh6xXN9k
w5Bj2XRNTF7AUWYx7SvzqjAKYjIxSG71MIBLjoQ329J3a6+HbMz+I/GwJTO+j/HwX/6w6+TMxp1g
OKwfb6y5cw7pZ7qcXdty0q4nh9QsWi8bjVE8Cxy/mbSi+/fWBDs4eP3FDHg/hW/i8K64luYbb3m2
rlNgsQWyMtCOb8WcZgnagfBxYbdPClKsb11RZ7IAIgaMfzTC+VOMH9+gp7r8UQr/V8dj7OWX7Fma
je9tILepBYp4ifrbOVbUMR+pKXhaGKHH54+O+p4fACXCLn6XwT1jWbbo9krA3GlBaQBpjjRaboC3
ElnHSRsNIL+J+dAQMCwtXjs+WHS6t3WhDdmVVH58FvubHIRta5rzgZd65dQ5YZVPH8Z4ZW7Wf23u
4qU+X2DVXrdmMKJv2AzR17taPCHUANmFumxtlX55iIyjd23q80UntH3Z73YSR0hmw5I5jFXS4Law
aBzemXgg25sMgn+O414659BWThKX2QFSfZZPS76NxjIQfsL3/YW/vXmG31oLSB/lcatwW8aBTrj2
PUq+wIhiAttymS95qcBWQ/73CH3eeQSNPlnsJJ67TZXeM8tA17SGnV7z/e460ZuKtTeeT+9fG6IM
LN9Oj5mg0s4PcJe3KtYxddwKWgoNjRG0Dlo/VIIj7GA/XpS5rcy/kb3Eej6wKDsohVajdB0Dwr9J
mu+JuvSa4bp3bn+EOl+Qnd8gV+gCMC4IFpvjXICXuru49YIJCdCkO5Y2icvGLKxr+DHXNs3LCW4r
xgBLpBeuL+sAon+Ix2am74LHqLAZcbXFk2xjlZaWDUfxKtE7cO3LISNfR+k79ahppqGsWR7lPvBI
GCWXLhsvpo9DE+F47PD1DgdjQnG6b/3fBFpeqSXJ588H6PUqbV8nj001RkK6rCqt6kivLPjD3hxh
4JOfux1s44qqDZOXProSazjdUmF6LeCXUeCya5/XaRTsoBUqJy6YuUOZjo1ILsxa/peS7fncYNgN
Sr8JjCBaktPLZCsbPQpiMDP2p2/q9kcM3d9PgsUmFkn/pUqUl5ODrUum4K5O+pbY8WF3SA4pkDtL
eNULbaynE/Cn+edE4WsVPe8qBsIG8uJwV/9IzCQlEv8niUv1eCtbY8U/V2rYl6Qq3/b+zwKpQpbk
lnWcQaxYz75An3Y0cA9ZkV6RLVKqPkT8LW3piA3ZiGqqBCdNQissmn9LT1NXFet/+ajayK2RQ3q0
6Z+inwk7yU2r481JlPdBYtfRCquQlCmXU/sjfRo8Czgt4/IO3H+TU+EaqNHmjNfKP7BeAXV2dLEt
kUZTbtznyhERqLSKuwpN+CrDswrWdoDA5rV+DccyjsvWuwL7KV8NJcGmcNuwLMmYKfHMUEwUL9Uz
hR8FnZtrRTkjOTU6UWOG7BahJbLRJFGETL4FO0QV557vg/LrB/KXxSryMhwIQt01yNC+Fr4eZfUH
iFu5qVnRqLERSxJ/nzzAiKmP8aJWz1ecp7NGaK7hlxOdP05JcNpi0tBPWVAMQt6Abp63Ffmm/vEY
EL1wttX3ADcjr14gJN9fuGFaOUTozPPftP7y2R1Wr8qG1u6qZJiBT1yskZX+pVuUaI7e8DIoV2VU
AW4GCwC21TpOI1W4CYwKpQ/BvMvslvNPFMcXVEd6Q0FQ72ve2c6LpfMPh3pY/CeH+ipgyP7nlImC
ECcXIss3GpMNlByM74fEz/mlQWW3Iv+GDaZmmKwsRyovNi9EiE6eOjgiZtuWfiJuda1C0IHcy8CR
YY662Uhs5zxzyAqH9pvX4yPEPSMOLUZ2LirkphxZmfP/d9hpTPZaVOsf8m0lbEV/FZzw6L/UV/3i
eO3GcpbU0bQgBJaFro6d2LxMxlTFjF3ardhfwOaiNovdo+9MQ6NYPg/j9SD40VbdYbRilaGGO0Kj
lSxw4D58ZlePxWvbd8No2fP7JMjgN62LfnfdY+B+e8Xl4hgIvUEeomi2jVZAXtpNDefivxH29fGm
dSZwj0LeW5mxJvKjvWtH3VCf5wSDLhuQoadXy6lgzwuVbgrq86DQxLbErIROOwTM3U/ETMb98nws
wQldvQoGrFzpn36t7IouytrL5XNhpsFgvKCknglYwOOjDS9iufmzH8JRWV13RRN55wzoNVlRpt80
uyAQSVBlNIUwae79Uu9LokJfryNvr+bPzrGLRZAnYBbw1Z+toLWuR2rOBqnA1TwLWxbG9d+65H2r
oFBJls70Iwgvl+vxn1zXqjpjhAIroZSngZU5wYktM8FDxLvnuwVJq0fXs9HRCYFx9bcR5V6VFWIM
fX7pSSBOkKLszoOBD0aW+WLs4xrRB3JhDuZLqXWOIbjXkx8GX18VscPZTbb7MgUCrQcY1FtrKHym
xYhqwGdU/3dSgep1ShyYacGgDjQv/djscpjZVYlz+PO+UhgA97Gu4SJciLNgkXdY/wWo6E8e7SQH
xdpiRcNOwNmLFeEmhKe2RccweDuOUY4pkHrSb/RUx1r8ynf8IAdbHKu2yVTeaPx4mVDQOF94ZnDp
gXTXlR1Do4e+VG/GVeU/g5ECTcbQc1BVLBaP1I8C1luIZoHDO22pRYaT1LADpzgWuuxpmCpDj26q
zke9/LXIJJpreV7/SsG7AUq79sf4pAxVxjBA/seYjI690V2IwrJWp1t7YklYQoWrQvRDSJ+Hfcyi
GfzJvUKXZWpU3OIO03OsBeDMe3m51czAq4Ode0VKXBsuHq3uS7shq1RFC0WRiUVJ66xMKjTQ38R/
LgQZflZveU5S4yVSYBBT+xK3ZradIZlKwAexf8XhNz8nRXV2M+tljCh/9pG+bAfmaYqP9gRzQJXG
vvibLOiShfJpsLWioBQUBWAEDbMZgOlTYXL1uLf6VF7SSwnuHBuX4dWtT0hReppd1piMN/0XbHn7
mCVhHyJb/gDp5CDALMeM8OVcQO05pjCMbjqL0Od9Oev9Ha3D1KLxxiSIabXGeva2M7sQ1+TleW0k
q0E9VWWcCsDOIRruIjto+7O6f0dW+xeqHuFhn6bC7YXLGN80JXTSiaLrn3HIt+XBf1FDER+TVrYu
QwdIwKSGsFQmRVXqFQeZ6ywOWS3MC7hvSQmjLOMQDilJGxgF1n019W7ZXBv2lHG5kE/7eJ71R5m8
4csiQaS+Bleze/QsjZAIS7iqhFxqlUtvyhf37Ct8W3piV9mDM6Pa3+/DJ0jgbjBatNWGT/4WZlrE
KrmOlU9qdcT/f7LYEC61YVZ3yX5f4yiOupldopEgrxQiIqjslU7ylOS5gmsjaoHA9ivopsHjVDKB
5DGO9OYj/Me5zgCZDVCOXOghvDFyDmELnymiMP7xW61MT+SmaDekf/3AfIzfim5fpB5ZtTw8UznJ
vlLFOsPBPeumexq2Yk0yLaqynWhqHESdyn/xDkvsxCtx28GReneH3M+YKf1dycsnqg2gZeuJphPI
706WPd/n7Xc6hl6F2PhfSpwvKt2xC45AbZcHYkPdk4rwSBYNM0Ux+Ow61vhyZXjbhG9FdQTfvfxI
f3+vVZVyD7XhXVU4I8JHSa9KzL4ikcsrzvGUXx+HZtpAh2praEm3oyOsrZdJbq/J2nUb4xECTcL3
gtoR3d9DxDsy6fsPxEdYhXAAOTcnYYRwdrGLTYSBdfI9utkPGj+YBvvOleeQk4oL4Q4PKxkF+Tri
Qi3DSlP+jec3rxW+HT5qDJ5T1dzb5kbKidtAk0u484+xuYmx6EtLAn5g2iqFAT4yfctUXB0GOScx
+uVMbw2c32xlC/WCgtsTJsfhEXeY+7NhhRrRUenLc1eHPPYET2WSrmR+OIrSBfD095E2pztdFnq6
eImZfsFroB8CZEvDrqFe6txvXKhebY+ZF69MyCjpUzFBzWNicd7QaxTBs8ER7lqpWeIn8mvQ4skg
GCzUrhIl5NPVImIYaYwZDDbJjAo2EHxPNkqMqwp7Ev96CF7+CV7AhBSuA68Rkjl8QWY82MKOmqLU
7bD4xWZptm3ysICvoaUShkFpoLOplEu9J96JKEm3wlX0jjcwJGUqXGt4vrsZmHdqyUZdw5znqx/B
yjHc+RLK3WsyUZwy3oJTci9FXoDUkoSri5MHobSOMhjrSi7ZMvVD9eQyzzg2wuvknrhVFTtUSc9U
9zZGgR3WiqKAHMBbJEpvbbDrHAKqRkYZDqVwiPvZ4IPNrzkq63KNtd7TWFJ5nDcFC/AAXIUe4DiU
zcn+JdfKF85M2NezBqn/UI0Su0bDVlXgo/SmrWj/RcjRa7YtF2osZXfiyXxzl3vp/dxKcoURE9QB
BPAi4Z+1c36YY7r0i4jsWGgWlqGkwsF57oasG5eMgYHtSs3W9OToujABcaRykfvTKaMSlU+eIoya
/XLT9nYU+BD8T7vFlCaWLFGHXkjqxSHoOcqGjT83hI/T8lGYi9fSeUdM1DdIL3SRsquDZBK58b7f
PssIuFkn54bCQaQOHCrmhnObrTTxcS25PYnmcTXnFH6qOQLDemA9HZVt/FMgiUWm6Fat5Fz+0cEQ
uSt4zNkNwsD5njlvatwOO2S+nsyHJyII1izNvCrio3BO2n+AxbdN5EjsdZT4cqHrB/d4t8eQTslj
XiJzSOuOcynwehfEXkLtPv8Zr1djTtBzNF8IVSh60f4RKbYEWcKAtFduIxt/ZWVMzTbgzVBMvZZB
pJ6njHSYp+gLhVECMUYGH5ztoKgkAMkfYxjwYxC8MbJpOcKMP8ARzDGCKWAnKYueo3uJYkKq9Mtx
cmEzy1p10rersPs3t/B3AiOyB3mR3bg6hVDrsQX/4AF6n71OIzGzNxaz1w8zdhoWDr5YZoqgHlYP
l+PFFY3hRK04NcS0wkfJkSlxq/u5wIgPgsoCwkizW1qSMjCLd/ktuiIcuxLF674imzwKN9roFgqY
8bDB0LD4lp56kG89CLQllDDvlnOcSKaH6iR0zLjts3Yfd1Gbr3DR/6qCB8/D94miHGI717+j+pR4
4K4wLv6a5VvqvVBZj5jvNpVk6rQ09X+PTmz77j6/ij5DCzTVEYsHlFWrNWEUx70oSYCGll+36oRA
obAyB1hberY42ukOjHbxpVK45QH9geokl7s6tWvNlV/Pz4vws+dONplCwy+88OQU5cZzB5c1qWW6
7HwjNs/ieSlBMcjmCsN2+xy3edptMm/PDE2GuyYT4ORx6xgtGnBqQ2VP0nuXMmZ+QBvX0f+AYCsT
IN25drXTlUZqcjYUkq4SGljgysYZX3kF9L7jP3ZMGok0yt2+n9jFgrBFcKQsxJ5k50+4bhx+b1sj
fyJMqxcdcO/Qr6epirbS4iAuFFZjaia7Rzlyq32txIpS3IQ39oItLj0GG+R6fAGu7vCoy6p7q3QY
BEdiw+N33PztUsm4PMZUKzbZWGTWD2sgDTN3r9K0gN0mvnhxFwZTZbxoyVLQ/RJA7jbxP3E7XYJS
gd4A0F8Xs/wzsncax6ys8OJjqve1DPIc+wg9ndz6oaULz0FfH9zseaF1j13dJykM3x+MpgBfsI1V
jkwFpl8G9ZQOzsaBN67V30p9mbkVgXSF62ooBtaHddDi1+ui8IJwW8mG4AQPMWIqu5CNoMxnMJZ1
IlIv/5LGkCKH+p8J+Z1eIYAFuFeBjD4UBIgzZER7zcyUgFewjAg3C5w3GCCYLM3s4OvToqQOs5oK
oCdiAuDmXFLrzqJv3/Uv1iEUtJCoyN6BfZnXqvqr+OowefHkWhiWr+D09CvO9peZ1IOkWrTaW+Fv
jjd53b5AXUtiUMQOYEPE/EoacWBbKa7d7KkM0sIOPASBLkoxSUxX0DbuOE/LvwGPYsGWV9aBxkP7
ChOs6euNnKEkSaoLCNVbVHy5Ys3c4AhXr1QZtdK+p6UmvXoLkZTTxAKFraIDuCrrZEcGAhlbgPLA
y7inuOQAWRbxVe9f01gb2NDJ5KWcZVZdHHYY+eBtdEj9rpqX6/e5gv9/vwnxGhFzWrzYuF5VUKHY
5HJD4Zvyito/guiUjaO5R/EIErvsMhujrG948F3/mco0e7kYvjlyvbTX6Ikzds1bx6FasjruGQwc
IPL/IwKxeq3OGFDdAKLP5imOr4BA82B0dEYuG3WEIg/VVfIkgJ9iq9HwoibEt1feUoohEIOX8mAf
D7GCzEqwylNcsy/DLiQ3JoZlYma+023WIQlE8WJDFZPBXoisaC8Xzt4hawp0QiNkSYvy2thDhLYR
jlWIWJcLu80UV/aAJRqIFI9MRKkebEDMJZZ0/Vy44mPlKGNqmNBb/u/WCg3Z8KHahtm2TipDf7Hg
hx1ByUyujZVO+dyxfxPEhVrrGhaIfB3mFiPR5n1Kuak62K7zH8ZMVqrVE4kpijMNjNrsL6Nk0SZn
mI3FJXRp+fELpeBuxCtyisGRUUtlJzu79ECEBJZvFyI3OMUkAUAWlWZ44ENHSW1lHZyRKcGf+DhU
B9OmDrUYvn+0245M/cxiuxcxjidyM/bL/ZW9HcAILOjFjaaqypTdPbBXlvbZxoNSS7vXfl6AV9cm
ukVIoQDqhzrbeiOZoLxOmzRYravJzojJ1XmXswSukWIVCSokvxdeG7W78PtcTwFHn0+knGoTM4OM
StguJKgxYPeqqL3wRFRqNdlPyE64dJQkXLzq5nSB3Iq7VOjpHZX+VMUikH7g95/30b7ydlcf1dKF
Dsup4BzR/wDMN237o8AJwEZ4X5TX95Epa0+YXB4aJuvAJZgDfHe38j9fGjlcxlQ0Y0bp7TuiUCQG
4mhi1K+4XTrjA1qU+nmOV+orXVE3WHpjIwreXKSl/G952Pny4kMrZAvPM1pJfKJ880+v7Urz8Fo2
FIdJNRWQrrpzzzqSaG/ECFhdj8bw+OInqh6oGgY6ngjObbxBabaFPIT0/lZgAHctYzaR2ybT5Ngq
Cf7bw8xK2U+paClbpEgTIvzebyyuk7cCEgwncewyN6G/vzIezwOawCL/wbYFXNGnr2NQE/eZYZcC
UhNQJ6oqsB0X21CmeClZZEE4rNN7BqNQVCQyMjDdg8DaLyIWo8izqhFF5blXr9YpSvwBc+gTQ1yx
u+2XMN6ctYSXsWibYQIdAcxEnkvp5USdzsA2VCz5LYoWN9yAnRJNRv5/6iqHIcndfG1k846QaJDf
8h1gvOPayYYX7hWQCnSWHn4FeZy5h4o1cJFggRvej4Ggh9ypo41aFepnMSAyNGLxtE5/Sz6rJYb3
rauq7oVgxqr0X9mHrb8WScyCGJU92QD0F54PffHpBpiEvknQLfhgZHHQIrvxQRHdlqF5ZK5FSwAj
McdrFY23r681Y96sWJnPyK7QGc6EzsrCSiWt1vtYQAmAz7kRLdsicPuP+ovlPgZNY5xxF+L+FTw/
UME1hqujABF9e1fxdP36JKovsl3IYKGn5QwSeWvASR37JExDO/7eUglizHLjhJfY1rZf4au0RLmV
r9ss/PaFwFAqhEyLAXYLN+iu/jTmcSdrRSRhCEFefaCMopypnO/hoHHGfK8OwTWc9YzNawYCNhDa
0ze9+YixbAjVU/AZoxeoq5vpp22mZoo9nkJ0Jocq98BuGo0nl3oawrzPpTGZvBpru7DeArsVe5LW
XVKhhQMJFq+6LVRPuIIWicRUpoDxQodcSUOAwPi/CGijbfVyfash/7X/0/LKoaaxEWCYQYVsBC+I
ftk4GoTQYdWunH8UMRVETczOXolzmb7Q+c/roFuTMO4FCJkZGR5q/e+HaD80IYmgJmhbYp1jfuE6
hqN2k4+MFP80zfLaEYtZYDd8lKUuhkupObdmNF+vbM0rJRRQ1TQvNOLUV5QtSCvzVB3jgJm28ibT
oavTEdOAVSKXlrS2CYggcUDlrRuKOPXifDkcxWqszuPeOgrHvRyCqSsK/+QwyC22kjJALxEbfPj/
MWzYBYwiwGGFE9r1AONi1cObKMiG6VsGdRVO7UdzVzF62DEeDOMY+QSnktz9Kk7PC8mgaSvg8cqj
pd6C60SyTyH6grNarWs2JILIohTekVwUhHgbhIHto0luBUIITR/P5ZU5TCQe2M60QsKXnESz8mGx
myEQiUqVYxYGSpl/+bEYsm/GoXsaYivtA2xpqrBoze5nUhPvpjqWYnL7nYLlczsxJCD/6ArggG7n
7TuNFbde4PMQ1eap64qPhneaz6M9YFpK3CyajjDFgTjNl3BnzpvTkeMUxWM7eT2aNgGPTytOCWae
c7pwmBVfzxjaSopVlzJIwLpCmN0Xmt3OMXKOmGmdAUObn5PGYv1T/QgLBI3jPPg3BM+DSVmJE28u
kcbBn0slPYxpJW+lJKRPBnDP5JRv+IKQwwHO8Jg4bPts8qNz7P4I7Zixc7pFp3zco6d7qlf4HemY
ln6AvnO3IwPlsUXZpUWO8kZ/0XtzyK7c1TRnlXWi9w1XOWJpetqTaOe5mjqeusmZ1UuH636eQjUL
oYLyClg4+NuSx8Lh3MXnctVXbW67LsWDTXcKGTAkyiHstVm0SkxVW7V7eUjUSkwnFEmxqleaxfYo
hDXJKMN9w7qwRBs8KaYI4iVkhRymQI44nczG+YkPOEH8SkQ8/Nc+D7txnWgjdY4JssSmZsyXwaQh
7WKKL4q7z/nESPxBSvCxxh11FIRn/Evw/8nu0+pZTvWnWgdffMoE/MUZ+RdMYyEXCYk9LA+R6U1p
1hRDVud22uURI561OGLrHkU1PeO/NkpYrKsJozr1Tty1LRs5Z7UJh3q5aS89n1gaCdgGc3YkM1uV
liDXxbl9GDtwRFSUUmHQYc2yUBZ2VkyXBFVHG7e22T45R/vtR6RqfwawDivN80waBtxN1gdX8wHm
Kjka1/IAY9B6+KIH6S4L1ucLIW3OIfb7Ph5Ft4Mt1iNbdH9wRHE7FQnPQQQyfZRdYUUaQoWZ5lyn
SR5LxwAD0xWkA3k55p8WyUYII8DPFbgf01pvqv2rYGybLZ0cHVih7TLAEtr6+8FhXC1XVJocS2/G
Ubk0tjJwJfSnWUPkfWb2nqTMpYaEvDg6JhnP2aUfpdKUagLIiVPj79q0OELjYN1srxwlXqxwkk+s
x2Zj0bDACxzeeBi257LGmiHHvOYPo70kEKwJqiK3hzatfpON3VYVm2iyk8bK4TZVaoT+pCfLKEv/
ASVKY5j02AXcsAhucGDER62lJa/LZUqOLvK6Jf+qlHLiAjabdbUZDYomZBnzt4iu89mkk+zbeL3l
c8p73eyQrK+VvplZxMwT/xlnWV1YjuGiV6tzsA1SdkJHghoxWWpGJsWwnHLi75Pdb85S1zCTsj5Y
owDza+u/71ib0crFErbCz/FEA6DJ3kZtXNH27hEIRCS/Z2FlEBJe0FbZutiJwpmXb/KcqhIg4Q7L
455QRuREWHBFBLZMQ498Z6a3fzQPXsp5Sz5kmACzlvwtlMiTC0K5HMDpZtgwbh+vAyGq+vHyHzXG
yu9wnmhQYwERuuLmdbwMUiTL9vmtrjSAwduknXILJ73EktcAmLyZkR3yjJLIYDop3S23wwx6QnJo
uXT3EQ1T6pGmHu5nZEjZrNgD77K6iFWgMn7vDeEfUaFoEFuiN+6aU3e/E97Sj63+AUFsfR5lQtIK
sssFIb0xKt8AFH6DeNwUUQqwsU77j3wEyDq7TFUxIRPSi6rT5qAPX8l8W7xJUrfgIphkCw7ZB/vm
wsnhJLgiRxxnKHmXNL/Y/p/1Y7iGbCTtWJMVx+fujxIFItLMX3yzV+uEo/oW5qP08SWmQxFt4C5r
DWrLNQtrlVAIBLUO6edRLs0wJotpYuCRYG36NUdznAbxTC7KFsZgX0TOtXaWWZGCcxI1PfNtHkV3
R90CWtIG/YC7YE3Mhar0qXmWidJsLFVTnDB+IVz5tEWUfY9TbhXIfUV3s5u2Ym0Mk/u/36vvH474
VDzo7KFpUPLuSpbmFMg9JqB5kXPmXn+8KYhrpg3CYwu9Z2wjDVLZUY4zuWDw7f/BnTF0lYFmd+hW
Bre7xNH1eBwC02jsVeOJ5ULTVqy9ckcAbXl4xzGOki710N60DUVSypE0r2iZIYXUe+DLkWPe7Ek3
G5JwVzFJ6XN8zPZ5g6fZZbgFewhRAHUuE4S+6UgBtK7tbI7ozY9e5+noZoYqHXC6JCjb6eQ30Wz4
rm+FkVGPVJXnws26GleivziAQ2POr9KiZxjxJ0A44w08uF6b5kz38EPFGUG4ikV1xNLYNGxmx1ON
BWhEZvJ8clzTlWyJ14cDRMAP43GB98sUx1nrXuvKRxD3xJ9nP7IRxPhiYqTvmgwLhJFTbg7aoR96
Oq7AYi1YyzP20qRDTgQlqzTdZSoQ0gN4tjrWHG0szZ5bEz7/meltpr+eGuNzF+JkCeNcZkslqP/r
KHM3A/Dgsi4tBWLkHYe2mQxhVnr7WVS+FPrfY6XadmrLyKyiXtg3GqvzUFTtMABzfaamNnHOyLyx
EN/dKHvktwFiyK3IHdvVB5ZQ735YcSSFMrfh3yXgED2d6N/QwWRkCjprHVUOqtiMXtm36px0lWWU
DM4MuAQ1WPpG8hH/u8iZQQ/SzCxDdIMS/QnUzUgSw7v3wuVI53B6uSrIsZ6bOwLnoV6xvVc7JeaR
4wrGzWu4rcFuQfWjRoB7yAG5rLbCiRSVAceBe5KdWlc/pmF7ZCaFM9UYuuMUkESil0jvhlQqxO3N
o5BADqgq5oa3gWOvhWTpxP3gzsy6pXf1/hdZ4qTPkX4SIlgY3hxp1tHYWW03rg6fmOst/M14qtvN
84OsbCWeTcSdqvx/9/RtMH+5jikY5iDr+dt0LEtDFYeYa82rXwQqxLdpR5N6GzfAclV82Z5uqZal
ollku/RWjKkz3jyRQFuHyQLAubJdUIpEzK6Du+BveJhx5hgIcX77i5kh81fmEbGM4gjKnf7PuJa/
8zhl/m0PEyc20xNWdSr49o3xRRvXDSWAnFxwoHATMxnXhXA9F4LkgAEzEmGSzUNFtDVcmiEXEISA
ytrvf3/2tZeiRS7LofK9+n/qjHQXfQg4QI6MThLnWSiHAro77BbNybWjLPQNPrLTbSlSQGl26SZ2
3tZKjzntdJQoQOhltwVKrLTdeeDDgxclhwBK7kP1GXD6SnzSnoAEZBe7Nzuz91tqI6Gavuo9rnrh
VG0k++r+QRDZ1D3Ur5WOrWbF5e87bV3PjTPzeHnq6lk9wJX2ag77c4wa5CsjxBoo0uPZye1V8eFF
B9Mvk7lFbFW8CsGAqOvhYw0rbqm4t8pP6+l8JVW8fcfHWptVHh+DwfFV+yNbMxHI1ecXZr0ZhnzS
UHZxQU0nNTqny3bpwYI3ggJMhKxYEXEc3KZP5MpFqsIrMrcPoeWHkMSJBCipyUR04FUnv2XnwXWy
vAU80ALuPJny5DJtff5lTj6mNF6nAqg1mpEioDX1RcCcr76XHlMiRRshIWgAdCP8iG92/kTjLHkb
dn57hUTjrCwMpIUbGXl+sssRGPrRzCqOWSJlZBeJuOHIMQGBVRQS5xoOtC3xpfeX+YQ9ntF7fNra
s6TezVIIJgmAIXBNcmZWazSxUx5zVUacAdnHsD6eZ98xqyMekrZUsDH46gYvl6vSPUz/LCileOWa
0lJa9d+XHJqnosuWdHO5tw0Hj6Bb1EfnBbB0XPt2iHo5k5PXNJGNTCfcKNsk64iUvHRsdP+dJnS9
9f1s71in/G+U5CmqCip2Xy5oKut4+pH+a20XtqptPQzGnZsevqPwtCCjTy9h4f11FkNrwLYGuL5i
k2ylwB3OOHrUeZpw3cIlOx43LSIgq+OKbH/iPAnWAtUizUyEAmRYleJ2OyeJwCUrzUnmAzlGh2tq
2lmEfWtsWkAJYEMH+Z2FhvyIAb+fGYEjTnfmqNvB5L9wF56zXsDp6E+GDkhRYFPQE8n+8oq24g7h
vKOFR0XmdXcDbo9MheZpf0nLM2gMGcY7wRQWSMKmbUnsUClQ+1nazyPfJnuhAM7MhygjdlW2e5yy
4+rDfPvGYwW7AzFbB2Vjl3D2+1EWLUKiExtkCHAHIXYy2UQnZi/oZaNADcXVrSR3fGQh2Wpb4HTn
8zMI59rO/oxU6fBFP/cOR561uSLB423EfuRM54vuxkou6MRmAFRPMZhYUsI6qKUJbOJ4mUmdceIy
hJXwkunpKIb1VfIG6DnXIXsekXU9kHP2nJN1xR1VK0QKH2ZWHBt0K7UCBdmACYMJwqAGEBaCqE1O
cOk35oiu5JQnTCUp98j3uzKGmEBk5VyIyyMJQHQepY8nKpoxDjlvH0oIq/XWOmLYu5jUHyoXGQDr
zaB7RrxnpNOc0Luam+6jRa8If5ivtU85oBBPj/a0Fssg0++MiT5fGMDJojjPXaMGOWjT0nCgRe9Z
05/38tlDoO0yrT2ZeQe98qeomLMj5cZpzTB2A4l0ubAXRgPeSujlLqmHq1IsMWP61vo/7tPRwn1o
/jGmf336rBMsE+TTUaD+OXJiOAkNy3Ty79RUyk80Khv4xBBYq7DTmOjF2WD/1Z3kVKC8e+ISYiBT
KTPuk/JQyJEpazQzrVZ5yLSRLMdghRQBdSxRV/zBgOvU+ku24zpy1bLYmxGqqW3hYhvBQhl/7LT0
RyU9BtTXXcnqplAvTW406RuNyxqitRjLJm+pYgL6xp8rW94pAh7OCIoUVE83vXvYUquHgq/+u7iI
BWyV9QfcppH2E958iZ0GCvMiSyIPhpQDVAcHh9gN54exuRp/gNM0nXnHQuZPuS362FkPdOAf2MwE
mBPCaxQxIEODs2pP9yH92Nyn5QHHfYqMfCKafJD4vOdS9KVFCKi8WoQkCqoBQyPB0Yop00meAt9I
HPALPc/BETWwFtvOSnAOs9/CjXbrtqNQ7W/xUC8aE4dJbo3e3J9/1+0NW459yM94mNGja2Puv3TP
MxTSVvsoPSKIcK0g5tRujE6rmy1jfvYE/jz9cERoFPIu0Pa0iDVd3x8YwplICKQnjHs2dajynkBK
tp8pl67Y5+Ajo+wxl2+y3swkdtguXrE3TwVMJ1ks6k/Gq8hqH+/2GhnkqUqDr4TBw4M6+2CXQ8EY
h/GU1BzMZeyN1LsU2paiY39vsRl36EH8NvQdh3S2OggmfmBa2fnlEUIDCwOgKV6dxvaZ98FiWn+H
aSMge+lDt1tyw6TiBZkkrkbNBcTO33LkvLseGMjZzQg7BtEM5eFK75Lfops+OM7rTIpYdAxiyfi3
Q9NWas77UTQDHOlC7J+hVIvM4RvuV+1PJqk8BiDAHkab3YYpqRtoFhesCCVo4nSjzuSbkcnX8UCK
aoNZWxKTuzDmPUoD2S1g17qefoVizexey186cAx87Ij9SCw33h+mhQX2a7Z0Y1NADW1XqKDIN6V9
3bpUVG8j27hgVW99R0k7BCSjlSGnLAKXQY24SY4cNIfIEpO8ldApr5io2lmwUM+qwMPVal+V4rlt
rTfRuZWlTn4DlnZ3JGhVwhyyfj7SUNlRMsb4hEej6b6vYoaEgTNLT0aUpSjODM5xk4zAmwtD1P1s
1/Ak8oeEGMFHOkLYeJeAUicElpWMQBuVYE0nxdmyrWNFFaxtx8qfg2biB6z2/P0oHQTsnp+JJaJg
sry1LW5OeLo+nKmWODqY2Zkfv6mNq05hrk4f2kZYZHobabENHp6+mnNHjqXjCYjwVnKRZkPxOhLi
wYaHFp9zZSNIU7Q5VviroyYkGcXZKRnrNcyL44DSVP5lTP45Al4m6TYElZS+/wFDRNEg9I99Y7/+
qr1J4x0UtMJB4XtAFTycuqy09Dz3do6j+1Gh+IxQOcDSsLfWBpvUyF4eVH5PmW5c8vddCVzqrU1U
h2OW8PmDCC/KJkhRA5F4Jtjm40cTfIwoOfs6B95EtuH+TsZiA+aoZC547X8Xsnjtwm3omZ/aQUl3
U+zXESvN4vRmVJYOE+ZRpOf3+eDBcW2aCJAUBEAItpeJlOQA9hCed6lbsB556u1lzUYOjH1xoYr2
GHkOCjvWiLFwOzDphhHKKUM2LCBUTunShQT60qVxOON3qdYm/chs8W8+MkxFWUOwNIiDsDwpNMK0
7DhITtyiQa3gwrMk4YFIf9XEa+9P/ljwL3zGW3aDkSkLQIFrCK82iUmEIRseBPAdeXyER/jF4s67
aoYtBV26Wd7TJgfVFPYgoMS2mWK0sqLFU71hrvBBx4nQaufDr/Cu7H25AYAwThZFpzYH/3AykPXm
16h6nSygkk1QrCJzyzWofA3u9ouuRd78//da+dCaEseZ3Z8r3hnYVsWjjwSALiB4uuFIaY5Xv5jt
8esnaonUkxCK+NOVyB8/SVDfBlaMw3WiknDOYV/QtgMVoRZGBaS1sA2dUqAnbr611Y8pIoLvTV4O
Zz4umpRpwIk54dEITdPwiNDBjPsqKmppnsWbK8s8C/pX/7Tm62g6QoZJZo1D1KXTAHHmweRDSCCE
8SNmsoozElkjsNoM9u0Adfgp/R2vJpjfRStyHEa0GZSpWusfz5MDRg5SAteGMC77SJZkmlpqDH4J
9lX82/dHR1ak7We0iVdgGMWMM2tjPi7DzVYQux7mqS7UdzpDul0HYO2uphd+AMWrfr+CbCEMD09R
mH6FM4pCQ29TgCle+W8eAAxLRxpgxy/nGP8xE03NJXpD1axtmJi77qpdV7WA9dwo3cHH8DI+x7jP
WPJCfK5321KEAM2Hadg8ALWmb1yvckpFn0x/CZJXc5jM9BcifKB04v0TlP+O4o6cbkSd+C18OqJd
ZLOnbsWU2f4ZoyP4UVXzthLBqtOaD1izFqasqxRXMV/xPjsd/KIcdLK3yuT8qY6c66l6y9BjFJ8h
ZaiCZzqGOCwd2+kUClktdG0r7FHPRsESGmwjCnxNgk+OP+x1a99cS3qoJYtdl3tDSRvGRd7KEdpU
T/zUh8AihW/zbUyPjiazvmpyC62EDKdyxAN92IhvKPkGBp74nKKgW6WTZ/rGg04kHi+McxKreB3O
PHP9AOcSnM2NzxEjnZ/efb3/f9xVPtNIviCul2KmbDM5R0KxiB5iL7ce0EqtVHApebVOoefVPV6o
amszbz9aOXRQ52QnjahOMFz42A8H06LnJ8IO+7+G9yYUhdwnfxXOfPEcEGlGG4W2sLvgTsc8H076
2thwSZCyKRtKYKZr0pG2PBKiSeKUkSa3Lp5jSKtFMD4W7oU/jhxS3Hly/4WpSAccbDPRbV2w9tHg
Eh7Jp+Jxv3TBSu4OErqgHgVefMlkQ/FDEu0hE31D4jZ+v78qeAyQke+ln3LWpjn8pBIVyjGr4jeT
1eQVY9f/4/gaJu+C1+qrHFSqUDaaegkljXJ9gM7olidv6aVqs28QHFQc34Jd9iUnjoDsw7G/bl9O
0M7hGcuGOkEcq7FRXowok2l4Mu1c7x0t9L0uJM59Oho/bRA6rJw8/8gtJPsPnRIl3wVoGSEjPpyg
iHIV/Vppvm/7599mqhVKm5TYgQBejd5QInUoXnXxqlUiHkOdzFeDWeal4Ks75gWzewP5gOBoSCx2
KiB2TXH+N3ARTkL4FEc7afMUvr7UKJLVlSyqbukNjaOsxwlQypjzw//JtbDlwNcTCAjXXKQJAMV1
8rfJvctF7cYxMwXIEwd48JeVM/SQ0oinPz4FbGdjhw7AVQkU4FXafsp3mcgtrs21E//YEQfW8rzp
kWgnNRMqneG7DecJISyybyfTd8IHLh9PA4FrL0yAsvULLITNFwRKFbaF9s5C0HxWY+f1qGR+CgXF
v05zfa5pCcYe/Z6yUnxRhifnud7hElHczrIeDZNHxjrCVCgfOwxakVrzGWOYbQd4U+pglWKcFSZW
BGQEQuX+5VASqLQl8yooF6u9Sy5sRenBdP0WHeWXo9W+M5+85jS7zgA0F819kmrk2WoCgx4Qf5g0
0chiJVlHHuCPcqfHuzvNYxrog4vGza/i9i8JSXLRoir271GS3wY3ZeHKMPxS+SL7yyT3eMgUpBeT
QH2KXAuilJmb/6IAEHsgHxN4u3tFbOx+b43p6V4PqsF+qzEmvIBb0m1ItgMnVCUbn2vUf1DJz7Zp
kJQDi0K94CGxNb7LGM4AwcX3JwicL0t7RcaN0GBSmUbJcTq3gGMJpD0/IF1uLMzWq8dDniBkTQtg
hCrbOP0Q9pi5zSdkDNgTbVs+Az6D2nObSxr0fwB0f5QccybQWyUdhcYuAzLBTSjikz8QspbHtwjU
XtC+TmhUrPe7sQPmzd0rQsAzu3moyx4aTX5PJ9LRXShLBsBxWF0Q2p9QcpzB95+c3nQEJ2dqb5lp
9ktR/bg7m76zq7UMhddALNeXWV7kCjfrs8oOOv+KSn6S/nT7sIC1+0VnUhg/orwoPQJIMZdDm1Ba
6hredy4dYWQbbhf6DbI2DXVsw4KqDBriylP16lRmkMhyJ9hZcBBrSWQqPnddjBiV6sHmhdrfoc2G
WdDXtU1Jjx8GLFRqqUxzs41rHp5BjlYLFphHYbtsbpKdA7CyEJ+A9QBXZpPKcMlohZvs/0KH+3mU
w8U/qG2tGXoykX8lcS3KPo9cR6pzXXrmCpg+n5V1ZtMQlVsUj8fkhcokjVECOWFelbp/ydrZMYlI
DacLryTi9O7tIFtf8YKuBpcspLkQm4GEQB7v/o4dxNfFI7tW+ZIgtlLWsrQelGIQa12pfuAuoVOr
7buUTAPjvybKtLmYtH7w9Ar/Bq7XqvMy5VhtaEe3xBI+KIF0NVvogihfhiC/9IAG49zdje4K2M+r
52RDUBjpjP61h+isXHCw+ybITkRMe0Py4N8g3ZbaE4usF7s2zkrBpMA4pctaAOa6ak/qlKBJicCr
Eo/i1yATZJryaQ2J140J/ziIjU3fR2SB7YrLxnuPmN9HunqdGvvAeoUvh+9NvniqpSD/tIkQ9ael
cZs9HJnT20uw4orb6OGocpgHcpceiw4+fA8kpHZ97MVZwQJVSz9offcAgyIMByIZ/w58tZsIPZ+r
VXDszb2oz5nQmUAEGdPW2JUcJqpUuLmSM3fRhUAWuEbxYrFHpx/Unoi4qUicD3tlz7vLJpMNBacm
gaaGEOQkBw8gJyQqBSKUeUdA3BcBvMSsCB35RvZNh8NqJDKAD0nyUeJWKF/+AuBft/itwUkD20LH
EMx/wZKUAILAr58cNTqE4gS5IAEQCt2cNvafh2oCgzFB9xkhhj8sITeMVDXXUSxVYtuv2+j0mwcg
R5QgX+/1adFvvhxTGODePgb0FNN4YHv7SFyEvEssXzV7nIrsqZo0zMyCZTuUIimnFpnyUw4gtEqF
DTUgN4Y+eB8abmZSY/mkxzOSiOSBkOEuK1+0Z7Np8EleAjVNKekDumocoJ9hNEzO7+zWaEHFzVPZ
UQbBHUzMSsl2hnLsKZYlBCQomux+A4G8QwDwGqlfGaKqCwOcIn5nwPpwP3vGM4iuip5wq91QM2Bz
CZkBc81au7CodMmGrZzFYxAs9iWPW+SeIt4UNYQ88DdlEovKRW5v+N+8qgnjjqs1dCuJrVjscUIN
f8Ek/SFcVj0uztIheJDsu7ntqhU75QYoYOcO+ECxhW2UvqFJS4zI05ocyqLe7YlzgUYOwqbnLxTl
CPOGlQ40J+FLHImptwW7YEvPEsNB9MoPe0PDdciaf6AL7fBhSzHNYT9PEDJv8iyLP29Gp5l2L3Rc
Kf3AKLJrwvvXbL7rzhJqmuBH9enKGLfFf6ZpxOYWcHtcHZ51TyyDKdvCL19JrdHYDH+UOTb838J3
KSN8CcJRkmDaMfcFaGkHwWDnrDqJaCjVBDghLIrpY1glwmcBFk09H1v/q3d1WwGspNJ1bfx2n+dt
jr4UfI9D9pIqkHJKKPi0OYPRa7qoSHOAMIkQ5Cvu8rjQnmEKunVN2PVaw9Rqz7L9qTSVxGQfobzk
xBmPmIDxPY76V00/+qzDkiCPDfbh+jsd5rFZD91qfftX/nIxtWZD70PzGbRqGEJIexTZ4aW3rlc7
oQJcA2MaOmSLXZCxprfPFLbWA1H1ql0ksb2OAjO7Gs8ZTmRf96rRNGx72/gvJukHxhI/e+AKtvsg
I9TVnI9ONd/oR1712GOuKLUKW9SvnqkQoIDRKQvrZ1V+nl0pnXa5TIHmjcpHwDyXzG+huwQO9OLR
hxoJoY10Kz9UPORDqegjOgL3uY5i38ln8l/JzkaDjEQ5b57VbthXjHth8SCpi5b13ZhMTVTYh+1g
c96RY7Slaf9eplZKwnW4iKaf4GZV3TeMdWXQIXo4vSV9AECEzyLqSyig1/fiy0xRSeiBfVQxI8sr
BNnoohz92Jn7O7144fliEwC//kRixyQDcrnwRiWw8Ba16r1iHQpE/MgLrTJbpLIPIsOplboeZVMK
t1Mb4V/UHKCFMXPzrd1UfSo97DLPhCd1TA3hn1lWSveJ59QTIy4W/lTUGZXlVWRW7D96YkMLjL1h
oh7T11zF3wJxgALsL7JPBH5NZY5EXmC0gj8dZW1fY5+qJIadXy/V1Q1A7TSlPOdjmUv1Zih+2aB/
G9efo3XfKmWLEd8/3j/e7J7FBEt4aM+n6Saf+fvCNeoN55srNd18o5OPtDfEt9CqycwAMVTVeulK
tYl91TDdHQTAwa7D1IqhxG0a99hKV3Dy+3mKFpQyDxEHzhiJIEDPEGGM6MH6xUUiIWfZgQ57jA2u
HCqJ6vv1txkzEWDTLzhCVwtBqFFWlub/P3SYG/BVP56j3cAFGGcCv/HqOhxQLbSxnyLOn75wcsln
hhn8p9S2GkF8KXVOarb/4RHaks8YUcMz0clyVrEhTieSYuS/2hGLUuzKJmVtAy+ZIF2cUxoEQmf2
x1BQQ4z49z+D9JL1i0ZYTNUhq31w00G/ykorI+w2JgAqQOE5Diruxh+yOn/z2F/NE5tOPWQeoPvC
MwVFNgqEFCVwdA62yJFAyA8KN8DoyZpNcPreCyLF+dPDt/T1b5pQeNyipscmv2RUPurxb3NoMfdb
iemo8PpYdK9InRt2bgsoN2sQMRJZL/+TpOmCLC4gzVT9NCexGdw/3yIsJPmcDmT1TUm0DXSv41P6
leuFMVKpdbDDljImG3KoF/oujFEEVpSPP/GivFqXKd6PzY1HKc/+kmy1qKnuMfBJSpuc1BXXFNIO
Ft1rIyPKV3xoUv7w1XDOAKJSheMe8OXeQrEzv1z/pmbqXAxMW54iG+YlAJXkeQZQu6P/yA4LJfT3
6ih9q5cGlW8PyqTU4R2P2AanqJBo5tKqUYqJyWPIY7/jTdooQQueHRVAHQ0c1swjZcb3aj/RlajP
ZKTY0AuoriwhZ1hm4jTzH4ItyadyvtM7B/cCvmcH50rcjYkrGALrSI302NK9g3pptOi5Hn0GLqJ0
cKmM6anYz5tVeCzP2sEQIVgyi+DYYQh/c7V5aTzaesT6qqD7SArvBPomVPG0XVKjcex0CW+stxxL
1Fk/HQkVzsYjg9KvIPenoDUoiULV3y/MBH4OLDe7NOC5G3QOggTBig8GbOgZoTfsXjNPtxujCic9
F7bMPcUbffwUIJRpCuXHYbYaftGAg8Z+FqwurP70oMD15AXTFwmhWsVzy+xomVaFwcdPVQlWL/6s
tbdq8e6oFUwmSVPLOEUwH5CmLTKPtk+TRdSFvnwwInzZltztg7me65mQd775JGx6F97Axsk8Mbez
Lfdbnn7oq0BGUanq8uRhY1kNXYv4RbGBAtM4KtGY9PQ0n23ocsPvpSYigHn+g56ShBYtOSTk2zZZ
hAu4ShYNL47bmVVmzt67sO+MFCnyt4Y3hwpGBajcnYl8ntT0m+XGb1OUP5mUnSCpQnZabE9UnjPL
B4kXC76TC/e+NYINMksIyIVFbrMEBAVtl2SXysm097QLRtw3cDTcxla08wJvFozaPTTmrLVA4uA5
B+dq7xzYN9/jJ5QgGrcseK3fmqI2+YMMW0aAMC0zHNbW6zTRCohjJAu1ino336KiSgPUkkA5rkEd
xxiDAvjLV4wVAqn+Ri5i7YXPunNbSwbJbhs+qs1uzC5Nyf/cZLwksHfLYJMZGrxUV2LjC71/AO1s
KiIUi/K8NqiD8CC45nVNzxnXKbSjpuPbkQW67kFbYN+yeV2yv7amqbNb24MDxS/g1A8WlRMvGRes
s5sF4eNT22LmMJjZLeGEfxkqFBVSHHQSLdj4JesAzFVOtF6jfQJskMOTg9eHq3nzOg+ZBFWpzGdu
gvImPuet6EDUo7Q4fpNU06GGS9HGODKv6m76XWiiYwdH5hp9gC0unYfVSr8hhhtkOtHcSjDG5EFq
1CQT2qdyl/Rs9vlr+/6Yxsy61+sPu2+mxYw1tOxhuRDKtJQRLjJOUSf6OvZqyO4uQeB5WuWNC7vC
2bDZ2McQElkb8sXQJDqVYlGMcB+Zq/e9ujr/ZmpjFAiMwXvk+uhlEerJ+vu2plLTrxyxgKbNtS5n
E35+C3UAqk2wRUtSf4hfXYTxwRAfpG5qAVULl+M3pSgmKpz0bWJO/lgwRWMQ9bcxGsjgW/3+ZQdD
ZZQ3UsKZv7U/lIjZ6g7g1o8aG+AEbw08eHQavgJq65y88jP41YkOyp6aHL0OtasDRvUxjc2wTKew
e7og4sbqoAVVIyrzrqgvmcaWeUrqdrfEn3O9kZKVpkGnt3K5eUATC2Pdp5Yc2LTIdpJik+dLmE/7
KlUP2ZU+qB+Da0jYgmtp6y0oGURAYoXxcCXnBYlVy9BK4qVzKjPCnf0S4tS/ODAF7jdVYjA4Qd1A
/OmNdHbD3VlIfX+vGKMZ9q/eBmYa2E60a7hLtv2CCxi8+pPuFiNXoanKQ2+/brmhVdxY+W1BbCyu
UHi0GpuglRctB8B5wqC0F2QQUvv8rORAqVcq61a059hkGLonet+S/aaUdR4LHc8nPY5FaYCKPZgw
Kq/tYR8kiVCmU2OyKFt24N7a8KMTl1oJ923OqSVVcuHe3HTyZPHaAYPrS+WcRWBSp67CQxa5sG0J
oVivtUTvuuZ+pzWDUqD0tivxluZEcYoncZX70avANQdZeSflljhKR2S0YG+KL9O/tLY4oWqIvtGP
S2W3+n7odF/dRGR+zcN4N17/vPFXZ4fO6U4gw2MJOcI6rw1Z2TRsxA2q2aW5qzY05B7uKBrhHxLh
PONwAFubTM/CqD9zutOKxleATXZqMyGsuW04kJqj4tXDtT104HYS8pAYHx/p8lfzkauEiQ+IOcmq
J6ArPqvePhIsVrUIEH6VKGEC6TJg6cyxoORf5ytuzur1qEI2ieqCaRSFqFpuJxhFlrXIWlgC+Gj3
F8hzNd3rhND9j6HcWuJNm8ThUnnBq9waLiw1jm+kqad8dG+6D3XygI+xcXYuMxBKnzPBkRpDvp5u
x7C224vlbsjx310LSPOWNQhDziK/Xoa0HSWQqk5OlRKeFWYOk8O657rUYUZPLFSSz8RXa7S9irm1
4ksL2RnJlOsQSIVrDVrAvdsCO/mymTi7Yv670A00CIdEUtNYJxO6cP0kRC5l+cRtdq/v2tSdbEoK
C8Hwy0FbCM/E6egc1YRnRPQRfK6SHcKvChitvb3fQnPvglpd44ARDrCRXrJph4/uvdcPLrX50Z5K
KbBwSkDECQM0sumrpU7mt4Oho6/yBUNheP2L0UUgyZ6VBgc9+mU/R4b46ctG/i+zGbwNfWaN45Qi
gYjmXBgAfyZU6pysPvY+tVt8R8kwmyAdpGz+VlbFWNF4k8dpkC8fPuwqYuKENkjR2nqcjIy/luLo
lVs+/pUSdl5HpMlrR4FYfyVocOCEYTY1i8I1d9xOcq/jY/o2yPu7uNzCCE89LJMb7cvw9JwSPuk5
bs6zzO11cV2p9M8eUPc9eHcw1adOvXF5Q0Uk0Ske8AWz4BwSxXEwTvHynJ64kyQdqFnnt5BOZ0jm
DH6MaeAYs+HV8agIhZ7JZT9hROg17uZbMdl4SKb/CpJIRq2gaI8Y2IPXafJmRyOozqGYdtJn2QAw
wWHRuEJzZAYT1jTXi6b0TVEHaj7bdiEZwV01G2z6XZ0pdOG7i5INuyisMwHjBeMQeZBOT4+VTzmR
/bVC1iPmKM8QB2KmcsC7T6vkZyC5wejJ3INlKaajWTVk3Pt+JLmqGmqpSjDcG2gjn6LcN2Tk5cQd
vywos8lywBLBlSse10VUV1m4ZdhcXzqojZQv3LcwSEylhpMS4NtpAbo8WCkbhCSJ9Hbrj+5X43No
NaI+dRofjSdsLtkCHy4I0Bn3VRVjm/RgDsVC3so2uHxXsFlZgS5jz8Yo5JMqdHImA547imSGLhcO
mlaBHQt0fQ7Uqh09BzmBa3EMcZP/xd2MhVfSpnNRiNN4N2pDlc0lDXX4uIBKkg7hmWHfh3MuW0X0
oXq8U5WeHFZr1o0ZYxo5lWE2Bd/iM1P7q0HopfW5G8gdbaqKcFmlzyheONKHUw2teqjD219DlCHY
KhFE3I5oAwGo2AHzmC4KDh2LDoc105bd2aa9mv5mKFd+LpD7QUPVcrp26E5AHpiIwRMN/fpQ9nG7
fcSBfzV0sKBeTYTaB/0dSUVfF8l9SOHkHoAbZSRc/NDdYoCJgioH9mbaxe2JpxPDglji6jun8oO6
Z++I2cvEwPIMGuzgDScHkg4MO6YpmDL+9qfmiS5BhY00Vm63HBdqAhPcUojx9REZafLEgoH/V9Ul
cJ8YIPonSFNmBya0wtzsgfPxDTbBzTYfmHtFs5a0zCAEuVW5MzswPrDz5v8Kbd6MDJsGKsjBfJ5i
GlzRa2kVjaz+mMy69m+dMq5BAgbR+UtPBBpNWb4QcxG0Liayr/D4xGv/FCRAxiyemWixFXLrrgSq
ataeJOV/bYZ3G0gN3fte95OBXLtkVHETyZRG6pyKM0BvS6p1b6ajPXZhFFKTowRv9M/X1ZGdLnIl
1vzjNOxwNbjxRRo97l6Aj/KYc4mKY0iLBr3N4rNsjVW9jsophldCZ/seKDVXhSbjG3/C41CbqqUU
LzQMjMlub7gE3Gnj9tkJqsfPj5TyUYSwjOnYEicQi2U7hZMbtJn+3XXAxfDJ358KGCaezdINmDgz
sbPCKWmegf+45fY3AdoOivtpRCtgsQM6yzY7X6m3f7AdYJBYvgeb7A7HqzqB9XqM6w/qEpy2iKAi
N/Q3mvfdR8o4vsESlUvMh6m+0WYY+qoIIYaUZoHAgEUCK3P5mk3BQUxbne3wnw4c8fDhHQuOYSUQ
sXKfCrhVT9sA/JBWwAYdEh2Hwb8KHymvfsyfzLUyP1kdIRNrh2AvlwUkHr43WDQB+OpMvprUiN3t
OTg3ET2BUQ7XuWjtgYc5Sa4aevtMUcXfrIavJ/88wnuoVhmvSnSa4oIrJw+qh5FJX07j1y6MdUvB
u6YHk0KYWJSKDfKflpPMNBrzhkPpaPMPaduWG0WCjcSCe+s9rebFO4q1gfOvLQDB4ChtMe4ByKYy
VXf4UtE9IJ4alcoLnES6lcu9JbT9zZaO1nQyf+VykZcxiEP8+whrPYqqW6GZfq3baEg5nD9pU2o6
AtwBpo/HF7UsCE4kgaTkaodYo/+jUj9IS9NoEj3baF/R3iSj+hoPAuXLLt6TOKmYPeW2lAGhD+ah
J6MPWqAcO/VBxo64WRyFpTJ1IlaSQDKGvW+pdHtZkjmGEPeIQn2yiZnA9SkhTIs6aOKzmGxJEdf8
o8caAcoRrg2lwHkokAlcDvmg40ab/78j2VRlbcZbmDMtbLBI+97koYq7bH9n/sPgtzWuOOfZhWtM
7kW6qCxvTQVlPIZGKXp/YkKRNaw+BIepp6Pbk/3hJUDWnjY3jaoUY8lw2tYb4Og6fcoQaRpKNPiv
EdWUFbxZXnF5Nfg9YpVZ7YfvY5l9j4IlyyynD9n2Da44S6Ci/01mMw/x378yMsikCp4++YvT9f7l
z8ibZzPWklfXJpGmcVcCfcST3uO93bNvkiA03+myexWUZ/dbCyUI9dgwHrUsCkWy2TDeeNmDKY7L
Sff2dYVhxvlf3NsoLqn2Q27SHWz5tAIjQibloXVEC9EsRFqICZsZGgLiDzQ/BS0HxZnOODdehmZv
qJOXCM2SkqtcBSCZP7HOm/Dti5hE/kagf3owiuyO9lpzPSBNE+U1hx5gd3dROGyW1QN+G3iLoKDg
DffXSmGgwVfBnBpPd9LJ/muIAXU/6z3XmUBcmdJ7eo2EQKugAi6hUF7QD5ClTmIXJzhEJ6NLZMSm
soIkCxc77I26yHksUCoo9zQejKECBTee/9evd7y3MRPwkwHObg5x8SgZ7BIwlHhoFDXLr71EscWj
x887POnLYejRz1WCwT/5AwT0G6wUKV0Wlqpfp/lWkBTsyQ9qTNzRFR9Fsl+uZqZT40SzPMRsRq4u
cjrYxgL+LDo3QnmzqZuQux1wWdYW6iIkFn+3TEs6JFy9GKFh5iXuCUXux1tS0CQRNHOJLHVF9GDf
9qi8aPYwHlcpEg+ESbZqL4N1O/hLce3u5Y0oHB5F6iqIOstnAFYtbPKM9R1KkkSne7FvA6FSSQoE
XfZzDKCcL9BDW18MNqkXZJ6gSMfmCXgRPzt+jmA7RJEUTMB6WuNoPIhdd/hU/UW96zpaMofDQm53
KMKPPlrgJoPQfeOiM4GhPzyEeFQekDQgXnPzxKiVK21yu6DrivXbS5UrlEXLdplOupQew6ONnc27
JqGs6/T+eoSMTOcy/mez2sKouNt3fLJNPEJzELYFJar7hs7srV8GONS5o5omPaRWUH+wFC4ZLhtb
kBR6Roprhp9M0O3J66MgEJAJr74k5VsDA3CCb0E4htYZo3hs9N9yBsFctzUk25Vfeu5kc7mFOEWK
BfcRtYeC6lNwEaO/WhDGV8qeDr453lyZmXP92I4wV4v8qpx4mLCfroe5zOE3q4RtRmZFOymAO3+U
4AA+TBARM3iAncboltwrMS2h00nZixxnkdFAvrWD+8Itz2c5e3yMK8UehUszgmjscQRWx11dWa6F
/HIVjzIBbshFXiGgQB9j3zS4VbuKrL+Rup1CJ86o8l3oT2aS4qda2Wf5fzPUcABescMIvLhAvOcB
T0AGtBTxFC96WpUlHfGC1JTYUV2ylOM7tkakXvV3962zcLQkemczAUcKsi3y+XXcWYmP51IIRzXa
JQAWtwNeosfOZfbH+iMpHzhhtUhVaYjhEWD9kGgZDY5QAIzqpnUSDADlr1i2rzX5eDbBQQktOIsk
ZBNkEh50ABzoNtVA8c7OxB+2PXyHdqOlr6tulsxwZC1T6uPp/Kh6PmHzC2Vmfoalt6nvOE6WaEdW
sB7kZG8BWWnJCof3jFd9OwZNArE3eTIV79N/Ir/ohT9/e8XPXP6iw//80m0BQCZRF0WXEOPqXR5o
WT54KI9x7paBhbVcY0hJcA8JcY3Ji6XyUpTBidl6KH4155dO30TZsMQFm97zEuQ4Q25PZCOcoNZf
O4AX8cARkg4CWEDcKeU47JqNhWmkqZhryPxyVsr4ZK/JqPnG6ZsYwfNe59r+0VIG0UFTtez/f2vk
9DV525NR6V3sYD1uJnYTfDqZErs0NBjtdf9mC9hg12oi6tNVxNX1XTrMyrQY5Z6T6B5EZsrKZCLz
mJGIjJrkIJktW/v1elDa5eQbLRzl1Q+7cag3HNYDnOpfIFlY2NidX0KDFp58V7oC6nHm270xMRlr
fF7GXlnakc2UZp8GeP2IsPZ9322YpGt9LkIZrN6uHdhIfBTr2AcWIn+x/iEYmbFtF7KXYcOi2Hrx
AYMLu0Cumvf1K78t71RvRzh1o90br3eTM8oCQL6mUDZDqFOswlZc77I6SxxJHOTKdiFYmW46eggI
4D48wu2nUOiGihW0sjMR9sNkb1p7Fe+IfguahbuQCqHEH7465IHnn8epxqUbIlwyzqw8bbbO39Xo
eTIy1HsOp9h01++X6kahHGQda/7tkQCm/P+eTNPeKg4EGpO+aub2td5srBAQiPX/W48XGZ6ESUxX
ZWc9lzD2K7amQevt3lQutyT2n6WE8+/ONWjozWZAykJKfUMH3+xjGHPlScYKJ/vWf+XJymXKz+cB
OvBgmpeWBxvidVoH1QDdAOzzFKSpPJ52hof4F2g5LcyRXWw5Gfhs4FU/Sl+2soOYbFf1qCTip95D
XH6B+x6Oqu2m8Vni2Uck27jKr5NxjD1G7GGC2Qb5TVTyUxgTZzdgpHIXHPpZhTKaeJiOiu7noP80
T61KCkKoJK7DBcaJPOpZeqBPmhO1FAmm4y3TBr1KULK//4/3IlxtpoDm31ls9r6J1W2pMxUUILG0
jITV6e+pNdTCHq+GCsFarvbL4zO8OIyembe01xpQuzh36u0ar77U8XXlM/9TAZcASfZA5nLu6h94
HCdPNrt4ojOPTrruwFL2uDABozjiapGCfIakSzsFHRdxDNzB++wctzcRIgIWIQDg0aS0eEYygtqQ
rU+cKNo4YACT6Qi32UnPHuMgv9RKvrjfEKEzWyzJ8NglRSJDgX9v44vAHSkqwdREhcyLO/l1vvBf
+pscw6CWNib2fYy5KORfKDwIHPDy4ryH2tJy1Gaa3S9QPxIvIDdvyH8QKH1pXVe/JOYcdTBc8B+x
zdTs2N0vqVwppZuiOCgS/JbGjy35WozIvFu8aeWs0mLw7NCpM1lmx64b1F37gIjEUY0M3qxdXHWM
DsBUN7/PiFJk6cISq9tfwuPGzJxmZY/IVXy9SAcDg2nPngqdhMTFPlRCnMND/NswYRXKJRv1yPWO
EGtxOTlaFo9J8dALhPRBxQGSmvsjQt0gPWATNXa+4FfbWdO2nrosYgC1PtUVXn4GtksBgzz178dv
qXRxRqSdiWP74fTAwaMk39kB3dzGrZWoNkA/LJ+akkOpCuctFUy5w781mSd+L/N/KwCOpLKdkktM
wTwJZKS3agSUY+Oq4ZUppTZYrYsc1E2TGC7FwUsK8AX3gR9tM7LhgZdqRcDOp6eYExqi47WiI+Ie
l7M2xChkPODn8BzgpNKPgNhHZSBLZZhiuvMtmLE+ZChO+g7EE3r+TwlT3M9Fultv7hZUcPVEKHY+
YEqaaj15oROE4svhPgZOWegJV1Wv7U5QG78NsfVt3DXGvvN5UCRwM53TRqWpFb8ysn7z9LXEWRhm
3XY7mWzTMqN7vsgAl0vIFLWRWMRUWq6AZrwh/CZNjqUaHzM8nb10fur/u6+xi8pzEYMyO58/Dtd/
A0h1KJSNDkNmnMqnh928ylWujKD5V3HtomY9IEoUuzLRZ+K58uaChJlzhQD8RUFR5WbATZDKI2YS
gS+DBPzwzBlc8xiDyrZ250XhLuS+71Zst+4cFbAZ1ORgrNr/wzDGjqNGIwBLuDj5xA7l0JSIgV/+
Pnj8BrmzDnpfzOsOqHlqEPVxUwJxmBqHYXfkSNFiDRZkffcqri41s2OuhhajV612vj+2aBVkJ6yc
ZiJjnRZ6u5EgyhogvXRTFbS2lFKOsac3+FvENNcNTAQqTt70ixgu+On/s6+nEMqa2SBFKf4CWzeu
eJIYiY6YDL4bpoUPhGTb6A5nzHUVkL25g+BMICogOCREGLzWP3ZRvpLO9xTDXtUm7D2SESLyaPSA
U+PaEF6EuubD2cGVoFMAry3+aKTzra0wqsS8NQwdpcgZ/AYipPzTNWG4FLFUmcgvoxB65QAG7qbt
mL0w1eLcKV1/ELxcYGYx3gwK64S+EMvDW1iPZVFy3ztvN26QORfynoLXdwlYlSN7okSFmSNkM9Mv
n/AnUDwugu/1tQdGaTSQOoEmnQIlmLCiqZAfZEt5iVS48N/sNC+FLHSbO2MrlznSwQ1uPB1Euofx
GiXqU4/3R8WDf+OleHhBsWrfeR/jNeChzj9p0OjbHCzP3HF45vuvgBbBkSNLLFkx6eq7XPd7iN2S
KRdkzwhsib+hdIthSpzAiVKX7Kw16IZmfSy2t4eAG9OfqCuwfl04Vs20NacfHv0yKG4smhF2RzmM
LDHmxC6vmK3ZazkKHO9Q2OC5iR1yDaiArKPlT4IpLztiUywdDJSP8T68BDwPJV4UaH07K86mZhsV
oIqgGamod5BLYY0EwvZlJ81aFztb2oyqSOVAXZiwp+BGqQH3k+BcNHxKOmA9Tc0Bqgod7adb1KMs
cBX68X3jq12j2aqLTOIIHSnX+psa88NUUKrAzROgQaV01C3XAf4pi61IzVOMXPPEaREmtfEXar1Z
bZK6nk+fzyheHLW2irRwSxAFXcoXxkaTBBUos22KOTLFi9nljgMLEone27NY6VyQWk/a6YGgQxbt
l72ThbwqsJqr5sd8It70bCZwmsbqHqshOMsOLt4lSP5LNdrVrxCHZDbrStaRgm5imD7mQS9/WnvM
nJJcikvwqk5KEOYg0/uHDpiaMBqDsDFSbQ8ItXDegIIAFreNf7sPXkijpHZBOYkGUfTtSprPU9nU
wz14Yu6R0mOMT8XMuswuLF7HbT9Fds4cdiBwebJSSxn/rq/ik6skNlzVTwfkQ9YVT4FJSn9UpPbK
kinLwNKfgeKA3ABzqhQ2AnODUyDtN9AsVMj6NqaaT+2WBSFo2nOj5sr6yac+DpZNP4E4wThYQbTs
3gTJd3FpB2PC50dxSeOg5/eTBX6+SeuyITrI+qY7HJLBYRw410ye/a39wv8zFQtkTxCK2CRtofJi
b+fc/omZcfVDAsouqqBlivjjKkidzwX5MhalTi7eLzTVn435Dl4ifcVl8DeItvVGqhc8f4PUMDBj
r0C2XasQb4MHyz7JI6W00f7Jl6mAYHvke6lzqhzAgYC9qxVpsJWizaRwVUdR2QSJA4l4ZSmtwj4i
usMTsthbd0xcWVDVoCQ3jl+kUG5Vf+jpZoQBb8l5p/mo4LBu0FIUQgBnZprIjqMlT4kigH5VXWWK
k/oSqWi0WhXrw5j65kUgNvCtZZ2M8agTUg85WDV+tmb33D+F8M14LIKYJpv8fYlDbIpNCepmqDdq
yrV7ey3DCzwWbySVIbvmq7kebXhCSmoT6/hgoE11OcnGEGqxewMVZcRg8DYp7jgnPVVwh4uu8CD1
zv2eHB0B4e9iA0Hwmo0osPN3XLKJLnbhsBH2P81Rj6DV9L6vo1AVln5T7E4nhtCaK4XHmFst55b/
Tp9J6KU51tBTdgZYCOyAG/Ak5GPLY36tSlROWX67/Ag8kh913kFaTL+8IK2WqVwFgJHC+rymcsc+
wFdFsSMxdu7VCyLAxJJqImKArpd2EARYbNzDzoYXbf30PxQ+ZBi2yhg/1VQ0tYHSAgdJD57cWWjU
+UUCkEt6TWOYIlKYKb87AsVuhHpwKge8eSAVGLLN/6T6A3sAUfS10pBdUli8onnsV3YVrmMr8vFg
qcIXFOlfghN5jAWs5pVWUsr3tTc4VoR3VQaJJZKNLZidLMq6BWh6EL7I5o7dkrRy2s90NhQTlTsH
dnLsNczGiMpbLjitXE+iYLVrylxmyMIqHZWOis76M1eDg6D8arYlWH7FUhmFavNu4T9sPBdMQc+3
vD2ffUtU9y99e4C/2CVn79CHc1VC2SaQuvayRPmhMDTpFIqeDPnuKne29A7Synl7N+SBdmKrQLXu
WYGbdi1ipBoF+4mjZrNciP25cuhDPhwWNV6pViqlkm3WaiKnb8bvOP2LaG2a6pA629pVdx0UOGhd
qca5w7y88zVv117PkzlYvckVVy/0MgS4yZV1WJOqv844seLkC4wtS1wMH6WR9ebf+eqJY7VOXdCw
pt/3FN6Hwn6Qjx2am8yyQLYT5zSynRc0/R+egvV1EZ20qHuWC7E2c+Rkwgy5sikHinxT1d6JKXQL
oElX3PueMzpsq9ViIk0NV8PINP2PA4vmPtF0I2bYDauj9g6j/QlN8yLVgOVFzCP4pnqht/9FbrHs
1TOHzWULVjP3qaOZG7yBg2LHM8ZwK+Zn2+FRUdSWbFWtIjwevgtBOyN4paEup8JxZZbUTkFb2W7j
1nziXcdAw/68oFQBXBtKwuJSSnehLZoOfmGeuR3hW/h3FAGgI9fQgr+wO7TWxsuIlxsuZIcEQaxj
ylYypDy7Q8v0gk2Jr6/EPvUVui9GWLfkK2L6aCO4j3Yau7Y1pppuRcveixozsVylW+p16nvp7xK3
9PKTRq+jD0VKVIbQNldPtaGqCSwtm3DCfSYwJ262a/1tn8NIToGUZSi+YqkNNWBeryD4tWd15N5R
G+bmOeUup3VjorG+hZCVGyRjEEd8ocbrzAhU+gAJLQPAGzbj2i8THg6XWF+ETnBRs7FZsQJrPnhE
m5DkUXAZRNb70AKGaKQkRN4lBiLHbIJFh6hAe8zCGcyd49WfUMiQweuEk8eHzYUKFi+1DrnvaILW
JS8mNW/njOp19p6rKbArmabKVrAOa4u22VtYE/FNm9eQvh6zvleg7JJzph7Hi4ObvlmqkI5wx8xj
e51f7hueBg1nTtEVbnvhh/Em3ZIr/UaLQxCHrjPM+ZdBlNZPAW+htNUVaovLL4QfpFxcEsmYvnMk
tpO2ER58sZ9ODrxbP+o+qYB6iAsRA91wn2ea/TAj+KJqIPnIvafvQbqj6eUdQKJocRzvjyZSDxcb
4exhvkbvZphEMXNAQ6vslxZ8h5MteWoPLUJQu/8o4v4qL1milQO+bXVIGuRRswoRra+kxW2csSkP
SdV1vykyLE/j0TcEWAIp7Ep3n1zV+LWT+PLU8qtQQcGjrMZb7F5sfkZqQhxC8MN5x02jOwXfLkjv
CA7nr0NlHU+xY4A9Au3onC56lWSTiHQp/zMtUeFj67E7CKHZqY6koKGUcj9nrnbzMqwvYe5Bf79S
fA7oPhHxghhBSXeOEYSopZ3JER/EQJF8RbO7D+086i2tqZjSBwAqmQLqqqWLU3CQqXzwVXJBD9s3
/FFxDPSHLcfQwR1oTQUjOW6FfJ8bqTiGI+Eh6srSzonNNjPxVpNgOx17vCTd86OYqmxkK17htpb5
2YjZ2E/YR9X7y32qJY0dICv8aKda3P9Q4ZODA8yhZJjOftlSc+1t6Vby5xoPfeWra5frFqS+duoE
dHQePoL8lfFWRLLizvwmur0EqjF3whkIgwzJgj8tFt4HP/IveWRARGAY9bVgBB+BGdnNBpPysFd0
a3H8QmZeAPwysewUY7/8nPs71jNyKTIqX9N/ulVkCEttMEGEaKi6PYmj+O3z1nF0GaMQ+LJx2ngr
fnSObFTW71JcPgID225uDNltZ2u5ENTpi9TbwOWfYiuUjF7t/fO1jtrs/QEs2PQzLdOIrLMKyuxY
b7HsL9gzJ8BPmLoi3sN4XQIaEh+NfQLdOq/sYEdjN8DLFtYNYYhYrIGYjlPX6SFyyAyF4UijhQjC
f3waxTv878GokdlLkfGrE1UgiEVqSwwFdwkJDlbCSONS6HxBg5rQdNBkPt4KupejSNhxWk3x9OPA
f7Q2EjvCcWWvsnbnEcW28y01/ie99pq85s2a9Z50wGV5E6ZqV7xuUU2ZCZuXrhF5qzlF0KA8z+Y2
PJfCGoWwr3jF1NS/P8J8uHP1odijfKs8KaD3pdG1V97w9wk7lA8qUJlcZnFCBHZNzxTMveWIxZd+
qM5+agNqsDR3tDstK+MinlVqbqXDyRpqbXXTKbU2kGj4x1KpL4Tjn91Pp/PdsNj0hh6bbhZIHSk5
YUT573pracjLH4u3TvFg2IBW5X98Spg0Puzz6uKMe13SrQ1BEVlKO+6NeKaJT8aB8tsLnTAkZAJg
yAKmvJaw3nDkMPTYo34A3wGHk7mP0IlMcf/iuMiJ9Wx+q4o3sMQLVvivcNTqw/5wVZjYFohA+reC
XczrJ2VLgvhkoCcrvZL3Zw9jMY9ycROd7loVDSZREtIrjacOG40yHGXvFI4u9KaoLURxccQ2peOs
uKDsvh6jSrLUYag07/uCxAeVONCdq8oGbpk7TDwDcHkIk+02NmGdYNqbEDOTlyRgZFPtpJQFCiTM
joXniO1W8k/zm2OXEQrgnulh5POfY6A6XUwOrOzfSM4aDqbs/8xOL6mSizjo2YNe4lLyyDkNt4Th
EtuIXDUSOECHpg8k7D/cNbvgeQZCNU/1k9aae3pFUQpwg72Ed3sxj/+Dasjp67XS+mbnnfxuvC4M
9NBGPhujbAyfnMJuyrw7+UDo4uXntmFOF0FgO2xcHmo/WN7lTFoe7OlUMbNKmR0bnvUIXdkq8+Cy
vKuXlAyBwcsXe4Gy6V1K3rxI0EJyKjbdzk2LFHBz7JYMZL/srbBWWFN5hzI1X4cW2YPVUVr2zQWd
QPPNQhtridyp7h9HGHNVBiK15K57S4OOq07EWK1bIXAVs0+rnEr5z491O872Sr/dUSLCZc49Rk0u
Qy6h4BbIvYKdsuk+qSqw45ZWeEpYZPrh1fl2fjFveL1XvB49czDzSW8uLn5umbvyYU2ClPnLTFtv
TwOZ5F6/TUiMAK9GKm4ontDFJecs7UduJPArv3GVzFL2/MO+qT6LHcJcAFRr/ClF64UfUAlAQ07E
UtwckbvOZru3WeQKvpyXwMs5iWOhdhfbUZjg+Dht/kAR/aMg/Lhr2bWfL23K1Km2/EthXXkMthec
vJ1GFzbl6ihUwpxUdNT5Tq/2ng4u3HDKY9DIox8NSvvSh8cNE+6muSvCQpvwvpDG5ZvkBe/P66Nk
WgEOAO3IRFcmlP4wNoV9xjsJFiFevX2PQHSbOkEPWhpZGkvs64Q5o4urWScc+MbfGiPRuD7Kexa4
xsZDCe5RfPblJHUcFN3T91hPwVAPlJOPO+n9MPlqZzw1n2f1Dy1XaPDvI6fYn66OVtrEuqWGfkVR
I52hq4AXR2k1slYplJU+BL9fel7k9dTI+TgqfouG8RUV5vDxFlIxXC69qVt2xV+4rNkur0/R9avO
5lev2kxxnqwxpzLW91UZgiq3a8kwiSFPOYL7q8xE5Rro/j1ij6b8Y2jNxR4QVhfZR1YD71vOnTO/
6hfMLlPZsIE8sgXyVr4EsCqHSYBGwk9g+pxwrWQC6B0E6khdRutR4tCpXgPN8PPXRB4msCGDVXVt
iLJee6ZaZdJKmWPiP6Kx7pKL1TtC3BW67gVb5oQtcaDLyLZhDdBuuoGIn5htW+K0U6c/6oAhy1dc
Z1ThGm9/atQtWbKwpjPHQDQAZypXdgnAsj3nAk/zpgwPi03rW+MH9GIoWqMI1dwZytStFUt8OZ0w
AqtVLYy47wtOSpqOSf+fpSs9yshRSyVe7H2xFqDo+h4u7ZgHiF8WlCn2h5PuGHJTObUO5pbfQtge
PlTV+h+bNKBoW+BmvmG0WN1gd38t9vbv72u0cVd3/dgGwpzueKNVoX+F+YnGpJQjfPhye+RqytFz
EqsDv9sJKDYEFs92+1a9maOKGrAaCC+viN+NXnXpls8YhWmKJmI4E0j0l/Fd0378B51PWttjk7U2
qqT8oue+oL4Np7+SvMaOHHs5qPPA8R5s2ceGxQ3swZjjokAa31ttrBrBL0RPJQrPKFzaAlAN1/wu
rbAaEkSCOVkEojPo2aJxd+AIB+OGaKJVp5HyddOmVe6Yfxa8GD7T1JEAolfiYdFrGlZLKthgpjGd
7Aq5JTnaFACGUHk202MPgxpLZcwsYbxK3i5VZ3rd8OTFccEEaaC8PHn/xZXEwupB5LzSjQ2Nic0H
KoM/3Kayych+dDLzfgWJO4FbJcpP20OQhTX+ulIB1xI/WaU/H4UU4h+5csuAyxhEEC07pIsaBkDG
wIplodoSy9PWAx8liuLwvY9mqXiIFyo8sBVtzz6bZgViqk7ry6exRll8u5NbO9NFQlllldI1Ad8J
xgn0cWzRiVmDjHHADbhelmQ5Iat5TqvWYOnMwCbHNzdaBt7ofneDcUu5s0ryl/BMybFxRpBJB8Jr
6HAw3hf1fJpmxDnP9m8MI9/g64H9p5gWdlS3NtNtjOTBIYLYODWwx56tlrfjd7ZNtU7qkVdBatwd
vkmNWXrNvUCymcQHye6aMJOysxeENZtPACy4HmCgd0Ud3KGWBEzoKVQSZNg7BGnbMwo2KqmjDFdb
z7j/3bGCErUTBfs8IwakAlCR22aOYDpp6epKJDsIZMPrJNqHqOrgVjysFxefpUpHlglrYp/fxoia
Pz7fI897TbBVjlaT2VUdGJ6/QhVt1XiljUnXEXIds329pW/qaA65/oElkoxZoAo4sFtE1ORVhHjY
O1V3jI6qRRMHYRXSi6r7q9GlVPp+BBKHArRibYu68gmckavHvgeMDRql/ZyKRl661UomWzn9sMHE
wc5SIVAiKhmkHnyx/K5/WQDLbZofeR0zxurQ49LL+Eb4rNuJ6I8CaBvOKlZZlTFAHgoNckqH6IUR
qzKLUQdCpHRDfbxEjuF51sGfcaHgW9RNs4moBc4jFtQN/IDlfanYiTpNEhGCki/z3QfF3acL9zA3
/DpYEf+ioZJHXEurenXdbHFQskDFUknvobfnO7YUpycA3bNnnDEwqtDefqwNI0/9xr2J4kypAyTU
o5Q46ej5RtLANxcXgrOMPA1AH5P8H6zVfQNlmzDCfuPntERWey4aMUgsjM4ae+HBh0WBrkq5Ym00
bjvMRXYc+G5zbiuZPr4gguA4T3z/zdWqXgL6NjvL/KT6XYJ1pqK7/Bd+ncUcSZax+I3MW7dIp99/
S2adIOCYxWvV2+9imb1BVTq0Rn5ygA22LBC5fn3xcR5W/NdP+UY/Xg0DW5MZDlqTTSf4VS1ZD4Ug
MH+7Vll3ZIj8lTRVYwxFkAXSfweY9W8uo9hIXwXH1qWJGIej9Ylh+Can+rXzw7Q/1Aw5Z24WSxlt
+Ad+FamTREEEFimp3IAb+IQ/IA1lx86udpBGYktEvt7sin7M3zE6ixfyvwwIDT8hllFlIOu01NTg
w/mjS48AugEaFDN9k9Xns+DuAm4WIqDMa9v6J8eX+TXkMx1193eG+qUfNTZDP7hLzExzF4M38mlS
OxjcLj83jk+RsxsL+kjqT8rNd+NGfXn5dEsokIlfbGBgBNebR1C97LD3dEalRk6wAYjlXEnzC+VQ
n2DepW99RbRes0GypwkBMnIA87DaIz8wJGS77wicw55PZ45RfIDUdcmiwRgSKwMQjATAuuCykMQu
MXhv8i/vBeI9M04Nkf2XV+R29M+YaL6BGg87vNb+sGbW02I+VPF/XArPQ9oaoHDTYojYFMMV2hN+
skrOql473UnqbJtUz1dEpke3J9NHFPn/ZhUkMRTyaq2wM84elD8CrKPgq6fJGiyFzidfM4tuhmcr
3nKHsAQUy2DGRW4/SmP1LupeZ5etG4/DWM1A8ELsRbaoyNj58+PMpnlHtXqDzIB8So1h0S3CxquP
WqZbR2N0oRREZzzEpfgLOyLIk3Xz1srvz+V1IK4Q0t5som+LV5JoMChePTSiwBIt3tPFpDqn8qlu
+7/ye8ae6a23nMPXw+uxgCHjt8V9xodTiuZSEPpO/57x9OC13ZghJUR0u8t6IP9e2iEVEjb0/wCi
GxR0fw2lYrUS4JBM/cKfyRzE3SwIMPt4lvFyAThEB9Vw2AIw4mEs4wGdSonUxPTZyoMuVBt5W5Ws
kPLjrKW1HFe9/wQ3DJc0qz3Z06FESoJe9U6eMzbqmfuBs91yryfWA83BwsY9U0NHLqlfn06tkGcU
4lUTWYQR833+K/lQQwYjKtjofHKjB2Yrq6gRoUK9hm5nJk8+eAk4I6R5kLSkbC6hU4jULqsmTVDK
U7CHYeNpq42j16pRtkANsL8zq9TonIR74c3ym7m6Au0F/g/C9Vpf1ijrIYFoeiBOupisrIFSbJTp
FgR/1wD7uB62vz93ObrWP4H/3Ui5BTuoxxR3LwIOiwihwaSEL0Zq2+o9+muE6jfbZhzF1Sf41q9g
kYhaAeNt6I8+VerruZ2eaGlP/u51qnJmzRiIGRWkoZ+J+qnz+t9DtCgWKKol+yVNMCTVPPBqIq3h
3dvEciiJEX1mLLX78cEsQwVpIcHYKE/iLWp6GlmweQEa1S1eGIn+Nt2c5ALXZUmFuLlnc4tJUpTw
WHWIHlYXEmgwuUcOdMCwbOPoeja6h0XQzNAY4lt6G1Qi1dpw73qOOC5jgZI/Pj6KokKKMt0e5GtP
6caH4QOT6538Hlvy+yQOMy3pAJgPUxTtRjM48bmdfgbl8YtTxkUD+D8vsD5YR7aCOOoEeEgBcl/R
RVgL2i5TpQZMXhQBM/BTvfaDqGxVWcN70xJ6rPchrHXuOJiFj4qc6GAFHbjponnfIEJo/gwEN4pI
3RzBXo38mDXtxNRCMiwY8hkQBoRUUpW7YFJclWHTUOaSEKVCf87o+agbLmgW7yoG6asm3bIoCpOr
lkSt3XiR4Hz7aAImnYDOkSqJc4qg+71FK/6U561OLVRymrOMNSWnpY7VM0DhcE2FlEOAoauxBcBc
+JCTcAvf2M47ftRgt9j5q4DNeVKKgi8+58H1px1dLMZS9ue+pf/vNXB7PKvoloU2hsFkY1thBK+V
ntZ0Sv7JD8rZ/WXTbluagoa840dS0LVWKp2u3+2ctXpo1WFaGo9cGBdM7EZ090OQSlYj2ACYqmSP
vlcgp4QE3SSVMm6Wff9GqOkNhCW1GnrevnAZz3kp0vatK+jsLCVfwCutkTFERe/tRVKU8B5HLKrw
dHoL9jP/31SlokqlLItw5Xvcg9xN0SCEgkFRp/ZzHiJCVAwgWe7A85ps8VpJZa1NNvWEPFPb8Feu
RkhfFk7nNZ11dp1eSQNR5r5oqUfhHUjij1kQJtNfC+InbWFe+cpM2CSQC2ilW7U6S26Blx8WrMs1
pdWSZEMFhnuxEC8GK1N1PXx0AKQfgc9OpEkGQ/rUgmW3grYlCBTSyU/pJz1SpXDqgTIVCLQwVrUO
8GLPKKYHD4CRV080kBZT0vtMr7g4lYE9tttP9xFfznowKWc25R46wk7Rkjf9xXdnd5CnqXZEX+3R
t7DbCkzJzohhtXcf1N7286cYj87cZMTrNC0fhQvQUKndmQWsiX9tupmVz401+4HzeeZGVAyiLJlM
UWE09VOaBpFUyYXUf70AgEzC4xwC5+Eoe1KEAiJm2AtCUvvZUpqnZ/dhLfjvaBnW/UoK3tY/87ax
ped48fo3ghY/9wWFi3rFwkEukol11+os550JX/RmBfX0s5rJI4eqrUz0cNSoKpMxxaDDWxaQjD/b
ztxUjAcbLgDOVUnVGJIJU8NEKdsby3c0LupATocG66Pi9XTvI989qxyjyws6gZMjPwOvH7upHNw9
LzRmZyb4OF4g8BuDROpu+LjnJAO1/fxkIJUkltzIFrRVPi+tcUW0uvxWIzDMtiupGLymbKxLMdb2
O5787W64tYoloN/IUskdRmkfk+w7tBn92uavfEtHAjY2mq0M8aFIEOSW4yEGb/F7WwYkL8OJcvTc
++SExYn2j/lYyQSRBjzuT6QkyAsBDvCzSy0aug345Czys8rUiiQyYIbKYW3PKJx37S+MGXeGPJUH
ZkmgyPkJ6ctfQ5C/H5GVyqhjpI5cKN9G6xm8qrEGqq8zRDzialwZaGQVm9EA9LAOTrPKtqDD+du2
SNrlipddFq4gzbtbGADkktf/yY5u6Y+tbkUW/R1YWws92R/SD4Zw7aH62ek2LB4v4WSo0dtVx4pj
pK0dLcBDZUupMrgI71Czab3gDq8NKK94n0Sjsm6KfMJ1sl1hDfnJybbTc54VbMd+ESJ5gGWXswb0
HOrJEUY0IS5qpiXPgQUcwoaspyXEGFowPhScW0GfSi78hkRjCogIlpRM1aZjJVbrTslOPRs/qK66
5vahFZmDF/1p+sYUqMcnENPzupsPUT7Uhr/EwuCA+EKjtZkjSOvIeZwPEH2ElbymdsYweGXx26ts
T3cUHdXARMArmjI25yfUbRO1MC39oE5wQopXR4u5EhRwnCAjTN7dXifmYamk7C5CITfowI0uEg1W
05kHmmB0SUIWviArtk+0PcJ7nscin7hDgpo954Tkgw5wgS+XmQSPEpyn+64MP1m+m+zyw5tE80vN
vErdZONjVCm4vWKGDiFnmIgokDOq8yMBO8XeRx99OYD5HMX5VmLBNvhh52CINUsS/NCX5cO5rkjN
J2RQVkKKtDwM7wuveNdunejdPJhsWsRMi5QHetuJEr9QsTl1eWadckWJ2Ec07o6siBKMqKQYo/0L
XBP6eNYmteBUP7ZvooxniZzgBPuB50Uy5xM1AlefFt4q/piAMZdbynJ/p5BYAyuoRKE1m1rtw6D6
peF+5Rsrukhykz2WHy+3YpnRW96+MwSNwnBS2DkD7/ZWjyvUI/MyRAE4basrlQCZMLOcLk6fhzBX
2WHesYVGFhrPwpsGVM8tuqe0PqiO7Q2clVI9+ckraOIyo0HgQSrxVeH6Y598ag4DrDrJoLZHTP8E
8zssJvMcOeAtFBxvZBlYRxup6kuM1pxec46U7cgf6oOky2T6y+jDiVJjG89B8WuWPoda9HwtMkt3
jMKDr0BXsXF1bgJ2k/M6FlAuKYQfmNOL+ybBEt/yLv8ii3ODH4Uw3mLtfRi5Jg/uuJUXRqV98h8t
8o9izXEVTScpWjgfJv9Np5mKfg3ngCqu8TgY5Ymwp5V1vOB5Jk0l2eYCgzFU+zzqmHcM3wP/PrAS
TMfRzvZxYAkMfCsqGQ4mbtcQDeyIyM7egW34KtMqotucpuw+H4Q0Q0KPhGE4CY8LDjkMXdi+7qLk
XWooi0Q1qUM8Dpeb9uHHt/fZN4RWc7Q39kheg6ICNROGXEl2lDOL7KmCRip+E6ZGS250dZYQaBdK
WYblIBqycWgPh9/OF+VUy5SctkslC+EAOrvcSQD6M/gMpd/wGUxRo3vYhgm/473M33RkwHlwzafG
DtU7qzgCDalQdj4rxOW0OkRm1Ix2jYUqyZm2/1UZE+TJxoLWIYS/Wsk5+CgSivS7+TWPGojdhG7E
v6ps01r0rzfhj1p1E64AIrciKfJqzePCuMphaR8YYiYJiDb4XLgDU5QDF0g5hl3y5m+KY51lkE2j
8zQh9OmOwNCOznsY8ew6OEdS70+UpmH/ZEAImIYmyem2SA5y2m9UiKHPDy9YJyzLpvKJd+igJ62I
ZWughF2Fb6QMgkzzv3DDQJipO+f8Dv0TBgwuuo3VkGLEdZLpbMuLSdEzKOs+ZaTNldq37n/y1Ik/
w51JD5jAAvh6nVnsynahbEevXzpjw+0+s7EEMyezncE9VqbRP2mv8oNOHfadWooYuCg0cT7WQyv7
SSi+OS4Fl7a8+vqaE4zf+3it/6Tia8q/kFHYjMWN9RlgYBPk8IR3QQ0skEXbQZ5Cn6jDxAc76S7a
lLfcf7H8dFGxW02XKn1oh+eweiLtxkvcQ7dxO37WO9EtGppmHo2o9svUPDsdYCPtwzPxbhE2jPCV
zM23OHh7isZt4iQ3bxIktU+UDZODup7Mu5xk7d0JMOHCAzclICzJjBlkcCG3atFvPGNCLOZO7PSH
wK4MDEJ5DGbV44uPUVZMT7mpNFNp6JSlDlSS6Av4Kl81swN8U87FMg/gFRt3IFZ6dYC2fAnI/ZIB
3yvlo0GtCxtqpOGHV/ph8EHLV9olq1dT5U9Jpd03lQM1jVICMU4+8V5R8nEGe1SwAcB9C/1N60kW
4ppikx1O2837JFjmh1Y39yw5TC08hoWd4tGg/u5ANGl7sO7SsofjQOJgVZbnOSTxG8SmMMPGMsrF
Zg4URoi5/PWAjgKoYnGOXfUVp6oQtM+DzBTPKLbsrOHpkRUJL5PJgmkKwndSQa/OCq1miZ/+SV3b
7truT1PLK1PPEpA2Y+TPXjrZPjsrkZXgyWfD97mpBR4mY08XYSbGKb454cQ+d9x9iKUagKk5Ifa0
OQJckGHbtLBJyWmzmM3JYIwYGkJ/msnX29L1fxmajOZ7B/VsxUp3Y7elUOBuj380AaI3VFYJ/05+
wFeU+igqq2m/jok26JJGrdtlbtWSgbiCOv3rL1XrVyv+47Af+Q/Sl351B9OONlUA3newImNVSkef
xPN2agZsFMlZefcukxw1toQdzsJEiJ6F2pKwGY3b7uYEYPS8QEsT2h8mG4a9Rf4Pye33L4+xpXt2
WOC3I/QaZBnXPUmip+jnakyEVOk2kX/4wesICPiZmrx7Lpn7qqSWbedzN6Hl67pqXTxYnI3mxhzm
ao8uDa0XrUj0F0Y3IY3aW5oGVtoNXxgddugvEE6S61qHcxYcJGHrvQ+QeGfUIsLdtzcJOJo8fGfo
T9Y0eBaMrMzcqYPXv/7h0Aiiyo5Hg3FByYotUExJ4TH7RpiZpJRhcMwPTO7VJ/CTE72NeIKvBowg
vtVgcPlr+QZ4BdHpH/2HPyKw6RDN/OO6QLWQupbWGpOmBxv7olGRqEGgWgPC6XCaQhQv5aoR7AOA
U/BvNlx3KFTuLaJsLQbKttSivs9R9NwBWgUP1i8UGSeLpgLVJiD4vd4PghVoKjGrBa1XnYuxwrJZ
O2xz+P3BQlT8ip7xUqQQxRKkYPfNufTJp78oj5smH8JM+q7fGXmpqHK3hUSrDKdddqXnpbscnNnj
fktb5xCaG4cngl0HWjBV85zhLknI5rw0+Ns0AFKU2HJO/cOyjjThLGHYXCQFiRZ0s4vEFetBWXBi
AeTvUqHQD47jPRxuxwPoECAUUmMNcHc/BTsfThc4FHdYFy3KgYpw+WLQvOVMOt9ed5RtyH1i8jn8
l0kK+TafW5qoRGvzDnZz+X++9DhFxAWUmhFyKa+B3S68K4XXBQ2odvj4o+a0kz0I9356tNc9CD/j
aw0hXwvIkD+maepfp0QEOhXGcZc/YaR9KTW8pyL4IKAx0GMY6NpR5diSj9UJjWeVNr6CTaHTPSXd
LJDg7arVDTHekKQXfVKvfGu4b432OU4Mj+d5oNDl1ivZ+bJOmxoZzg5zkFVGKTxJPVc60B0Uaj8w
aR3Uk1mfiyeRhLTGK+f5vXwKakpYGohwKoY9bljJZQPVchwePOs7vwY2//Xm28Hs0CETM3lhNcS6
ctnEhTp379MO5YyvVal617HMiFKmi36Rk9jLJSiU3a+nhw9ZUnL1YvSDGGx84R9S4ihXRQa80Ze5
m2xcURP1stU83UmLE8jiukxw/8LcUsPJrmQ5Yk3gzmZjAu5ROcgg7LJKu5onT0aaM/7K9Jql2oGn
xKLPA347s85I80zrjYzGX10pQxA+/y3N1z3A7+mbadHHQWbsWIDvAjZ0pdRvDTZlgq+xtj1Nb6b2
+KRCFyi17BErToxDZlbLo2J2U8lv4PMH2N16Od5VB/dvzwE0ogiDEw7GsTVmsMCmy8aBHqX6u4vc
YMg+Xy7KfoNBWGP7loa7V6XRQQMaC5C7wqjeJmUKgopRMa4pCMjFc4Z+DTNHCjJXeGLf4oFklp4O
btLWmVdSXnepiHh/uv94OH1gNzFoAxUnk6ttByXH7yIbfzB6KP5rObuJY6i//vKT6ZyaBrfDUIV2
sRoNJSb657XCbffYesYDpRbtTsavAH/LLL0GnrtRi42cd5k08qU4D/abD1k7N4yowil8AM3VQA0U
v9Ao3xOMCu3ecCDDPhKerN9OdU4L1O0m472bqc2gLoFg44ldV0nJXTdjvgNKFh7MgzcGBbum5I9b
qDdGImXOhv1BgU4iHgSMzS1ui5x7glMlSKXERlDT/Tk+wALC+O/7q6MsaPH4ftSXrf3OCCMxfF8t
ltUzmVrJFUkTbWDkOADIJ8D8OcSpRg6VCVAweOGl21xUpuuIBULTNUL+nnME0CcWc9rdYdIepziV
4MpDPQRpD7+OM/b4YZ9m9y3b8Z5rtHHgQmYydr3n/7j+zWQ9LycC2NSNRJmaVlTDKzQehHO7w9dh
u1fuUeCsxFAZHNjja6aVGZwKgAIeyVbVr0c3jxhbz3tx/XDXcP/jexmntGI4sLyUKR6RtpPI9wQk
Oodbw/W9Q7sBysOtHl9ZS4I7UeuVK7Oxi19QyjPzH8bS/eDS8L9hUHQi4j1pzmaYa6g6OOea6OEN
k0K56Oh/qJfJveNDhjgfZI7sV5LJdK4RfxgXzaz9E8l4FB/4o2HRyIHPsu2UgzKrS/k2H+EJHzTv
pJ9J6FEbT/xligO2lYhyrc6emudCWDtvVW7LNKMbbjUMLXkmkUe45CTY3IksH0q094BUO0WVYiL8
wLO0U2NASjpVvFS3IBq0IBkwb9AR8+JO0zHQC8sJTGosB9JkRNMrCfgWfqapuCYIOrjuJqAKHW5z
JRM8XwOG/sSeZiW8hDJMtj2oVmfXM/EY6s86ppfBROY/GO1OjdXaIjtNTTFqGv0Hjx7Xk0vZeEUd
SC0xOavRKbMnbGcjK0a5b9U8TJrTHIZU7uz4FMaan5nhExaWz7XYu1FghceRcOo0Z57fIZdD6ZcR
guWVGipudzQsJBq6zkD+ZcGkRNgayzD3oFC6ABPHoFhWGauBIT2Gk6GA24fVCxg3TRC2WF3Kx+Ak
dNN+06f438F1O25qsAU4xd+rneh7uldp0+kothz4vQoWblly0Kbk8izA+VDb4aj4WbGrSBT6qer3
DZgYcb3UwN8rP4iJNQETnSKuuACQZuPzKJ/By4khS4qVfqYnIB2jKKIFdzAC+UaqGPYmDxPmRXT+
97/UqY/eOfaoPLJbmAH895qk+Aqf+Gc1UX1ruHXHa8TWz5lEqu6FmLrZVCmxNITw8PbWdIrlKBpb
WuTdw3aLBLdepHNiHnr/B5QVKcWN58OIN34QNT0Gm4XLl2t30tAVRM3WkHLjdxSU2XmgTVKRP/+D
p9SEby9MJIP4cL5uDml77kn9mvyzWYT0Pks5Bh7e8xM9v7rpwPWjD2Uj4pZr6dmPzXFGOrSLh6ZR
0/TaQAjweRp5mqomekkKhxPzrsNVuV3fCq9nrIKtb+an9bYrrMdxwNMDHAJ6njLOWm2zIBUmqSsK
pWAn3gCBXhBz51T5ORrug+AB+reci0sjLkzMU7Y9dP5IMVdboiph7wJGIM+7r3PZo5Sf39u3yjfk
em1LrNJJLaUVKqKvmuaq9QDogTAtS7fJ0QK6/3DA0zx2CrzGZSnPUGUUN4BO8PpAi1g60jq1RR+A
kxlPaMkw5LRC0d5wquhwYL5mt0wmdvc0FmXkRktqvEHNa9Auwht/AcBC+EC+frWL/2in1L5gYfU4
VZbB1NitOJ1mCN4Wum1rLb810Rk0vONORw1V+kE71YVUaA8rkML+4MkkvKAgC1XFc6Xag1NvjCMB
H5UA0fuMfvZS0mj5sx3l9hytDXpX5zP0QxKSEpAe18rIAzgqyCTz6qA/3mgzzh4f4q9nd2nJ71Xj
nmTnl/Q1NBhy399GQwT1QpsrQPyGEc90W7rNA3vm1ZKBMvhNwBxip+NPk4XtkrT4Gic7PlsEiGFE
6/24y4gyvV3f1+PJy0K4UXEWC1O4+7CcHQG2bltQaQAsNak0p+n01TqYDrkL7EVZtnXNPho/MQ06
XH5HH0qaeuVEqoEQd4+vi6UaOq/ExhmC+FylavHC2LMwrD/TC5gYSVpbNAZ2GQfE7snijVBv55vo
S54Ol6iFibRy/rQlVMCec3qWFXCzlSQHyKPTgMxLeVeBzQTrlYRcoVyNVybBsB9n5YrdLJywbEjA
XeDZv0ErBVGjHS2uGbLa4FtD5idV9mldUyixWPmCYZPymlVvxguju/pKe90zyr3SOzJInLmX7mSV
TPxG0lAfTGv768ymfz8QXyxnTTno9dF/EnLa566r4T/1H3gVph83sNDKQsjSM4QNCxAX1Pv017t1
mdqJbqwqbN+OKr9bGGNquTZy81L9WpTndgHapGuuutqaw82ehyKDo4WYTba2/aMh4+HAVsqipak6
QYdrhVQWOfEV8sa7pkRm3gVUOAnpUAg6nEYreUKsYG1Pgq9myvLo93uMkLMtRKBUNBNdQehfz/xB
D4R5XOc3QUk66tsPfZW3WhyBofG+zBqerM/Hjyni2WHAZOnd63J3Wdu++GriJ9TK980mmjjMynwJ
H3MNjuQVaTZwF/oMmqfog5NBNIG/OxNGFsA03Qx5ApR62oRa3SsaHVajTtkVIKHMbj6SVQRDJuDe
CZKg8snoJuhSS7PC4inzC8kXVabeUBXxO5ud1VIKeSLS673aPxpMqWX4Fol5yA8wgeTEXUhrGb00
JPFFpYWOXBcoaXJY6FpSN/J1wmyPojAapGD7a87revcbhhCUno+5TFA6CAvGAXoSkC5ZSAKwmZNO
K4Ip4UX+jMTlVAbogpVHWedrWi0PhXcO6ZhuWhuUT9ISLw/mVecbwaT8bbbFahtxz5psOp+UvQOr
T3LiUKCwIx5Ig0kQPQ5PDyHqlQr62tfjsVDuP7T3fpfwNPvz55qO7Q02lCi8xeDOMXeoNFo11VMn
uh41/P2HRLF64vJWydm0lbKoUttGyrIDIAwPXC3ZqkE6A6FXIRHDZybaSy7r5wmp0WVEVJBHB8qG
h54GX5pBGvKA2tBK2ZugtooBDPU0JNpcm+Vrnq6H37VQlpshpwsq0/m6KwSrtDub1OAg9wLpGqsw
Tr1CFzzbf6d4ULBvhuKbJYfPY/c6w47t1KRaJWU5OxChiPootPMWpxsFRJZLpfN/JvuDZJMVjpAB
dtyUDBsOBw7eJWMwI0yYlqv1FODz/HL0HvsewKqM5fs/pSd2b7cL+5kx8TojyDbIi16IsQDk4ILF
Vcf11vMWLByi6H8YmFeTPm1gBMb78J4Rl+HnzYHkSoKBT4JrtHIl/e96BBhnCDgEq3GiUtNW95t3
5q5fFT9aDZlXUgVjJ2PCqHuwAjA81ho9sDAdcBHqCb3OehVk4/YXJ3NaAfh/luLj6zvX7/CV21wt
ckwOtNO9BB50NhNx+7NH9BuNCiqSIxv24C2ZuSrkyk3yx5BkT5sGJcDa/liGPmPTlxT0K+TLj23I
HcKNBGYAQoVEFz5+ZKCGFfPH0nEbk6kwgoBxwfoAOGu0FZaZTJ8K3qAeY4tdnx0KlOxVuoFAJuDi
kQ0VdHCO5oRrxcVUFkmsAit6izPp3mZjNmnKPIsVG9byYewVyp4gLFNKFCSj7RlfJyi07krTeu6s
6OBxd6iNYeOEJp/TwcsoXSoUjVrGwY9gffcWxtigOm079/UTMSRtDrrTQEAythb3pvkkWiHB8djP
D7C0l8OivoWIgdRRpeldE+Ma8ZmWRMei8mFy8/iWsUYONKL7u7uu9lAI0wvWSPjyK4BdHgx/d2TW
C0xY7uGW9sS1FP2DDYldtPKrAhm5KcBXKBDrGVRzDl0HANVW9ye8+LtDKY8yzXpsSDm8/kRQwKtN
4NR3JzWtav9GRb8vSIrPZOs/6wc2BUOBKgFyI7ffJ/tve1qs4JEd9wksVCYOZTd/KI+9wdgHMCUr
w+3gG0ggouwyzPvxgZCvf1ZxMYyelw6rNpWUolgu5nz+NsjIpS+RFLjQK0rn/d1dG7BNaDoMI59d
4DUty775gwJ2M8hPABxoHm/zj0niR4LMfk0kfnjmvbw+bAZvGoJIBBFAZrfb9JO+RmpjcGltsLwm
S/yOCwXtrYVWZ1u3v/MGA+Kbs2y7nMBQMHuCzv/HhiUIK+4DzmfwfF/wedrZtugrR4luzOs/vG42
VCJjCMwMV01/V2mc8AWgkKsMuex0mPm5jjO+RMX9WttSEhqw5F1kFOxE3jUXiM8HCTFYQB8msyNH
ItD6GXQUAHgZsL+xo2IfRTJvZoKaJiQmrfn4FOUGv57KxkOB68n/iQ9dwlNP71FGKBRmfB5Ku2zT
klFDbymUSAIRjeU/x+cUEivJPqCL0Ld1OQenDiqVdoe1J07UbkPJKXWPAAggTnqMAo/dHjzKqeGh
hUewy8vTmuxHBUba4CrnA/VJY2ZiVk6Ob0A2X7XwXKGR2VQIpTv5NXO62WgkU9O046KnsNqIhfG7
rnCTAeQa58WZwyJXreFYlBzJBnckDux8ULYHUEpbK2yKGLUEaXjDCQyuahMydLju5hjAPOlSaoHc
vpAcBr1D3iO6Gtg8pc97AK7HhUuit0V8CPKp3H/ksuwcrjOj3PZ+jX7/uBFeCmXZRO9iiQX3SX7l
rPHQ7251Kb3HI4/7RD+G8rrNbe4Cp5fkvTj76JPlP4pYz5kmV39j3egjWEyXgEBj7Mb9AYpY7olI
PStwZ5SOxIP7U/4FNv18I77sgOmOHH353s3CiNUQ9w/eIkhClOqyg2ogn3feInkDSfzrvMeLWQJ7
XN8Rdc7cNQGXo5IpjdmStPFk5urJ/Ox6ZsMysRKVYPJSYcvTIfvvGbiSnkuWIAzuMa8CrgmxTehw
TmkfqZBIHVuYxt/JaZpWormr37djxzQr0mthadBmIGD2pW05b70Y2EPvz/vpPbADL9e67b3wtQx8
J7dTfArhz8d5XreEBRmSQar6G4sJc0NEjIURRpLoQDM87FhNhghrzVVk/y1r6aBvcaDL/FlqO0cM
d51AgvPuAcPLYtZGoLtHH8g4QqWQwB3LpjSsmyliSMpwswdglItHlEoMlvZHb47k6vq6y6aJJqF2
aSe6lPVxtRkGluT+2Bgvnq5YBA/4+TA6/vx8TnS76ZO56RH423jT+sAFjSo9QMav3pZ/+Ox8kCTJ
w1Bvw9AbWEUYuZeZexylVz97bmDiRuySpvPYaDM+e9kKqncrGkxCic8Fxkw/2bP94KR4Gp6LLXKG
Bi4m+Bs8bVwi+o1yKAtwmbho4d/irLSEnBpfvctNWc3w+hK+DcogTmSZ4HS2GQk806e5ykBkXA9H
NH3SQB40uPfVojHNBnFOlYvmqisBjeBz46/QBGauW5gXJ1E6nGvIT188PvJ+EgRuBoVd+RWw/ZYs
j3VzdzrofvHwIx8P/87cLzuObFk8PEk06YXb5RE/xZl+GG30UNOGI4TJVNanQTUP3Ng8uyYnt3ZV
oItuJ2tMEzh5ttxgZlxiOSeSJGJEyEQw84yum39w6uZMF1qAaueBaQAEoZ6t/zGZWV7HxPOaLAO+
e2qf/XmvLo0uQ0EmLH7wplWRI8foeT62rztoWGnDtHDyF3rawD/aZvm516kM1ZxcGVNJBWgCWj5B
pEjQFefh6PUbXlXwyI+aW6jERuQFna7BWsGmDkgkm+nubQSDjf10vBhLA+Lv2ha8mV3CU5Ojp4T6
hDxaMB7Jx2j+IkdDREHCB8BX9UaizNzaXse+GW+jcCNWLDmKH5Rq3LEiENRTfBYtY7Bb/WcScc4c
gNNAlEkeo9rCcf60HKeHtIxb3hJbWJuhl8GGXfbtDNZkams91ECiO5WlDdEtRZPUIquyckJfqYWf
KO+5vpb11zECA5NO/z0Z56Mwpp8oInlQTfwrYsb7hdbKEANAoHgexz0NRRANf1foI1ON6fKgQasx
lChEHlsKU7kP+augz69n739To4C5SrIIXown8gxkY5AEWsTywEG7gKlc20mMiwXTvo8lXRzwc6xm
d6Nx6U8sZxEAX06lwGOXqQBXsmNLv3N8f7U/2P3Ln5WlyY4Be2yqpciKJAIuA5t43AS4lrNwQ6Ok
TCcUSy+QDL3l8LOd4otI1CiiIzfObWN+E73ZSwGWxh5jW2LtUhuucF7VRX7Nj8G0CzERsHs9CqQB
AqLifJSHJ20RfkrTX7RXFmbMx71HBGg6ioz7L1FQ0LqyowpCKVGfRpEJTdjvThFixmPOrxYNr8po
pMqhM2wNdlnh8DB04PwLvjmIMSj5nnmBcmob1erJ6bNqVzrXB5prbtm35I2sKDCMjhhOI42mQIn+
YYtqMvbMqNxFz1fU5z9tuwLzoASwDVv3a58yWB8B4q7jIyBMDHVZWGRJYpJr37taclEznUulmyFd
q64/527r/H63FSJRAabGo9PAMJYyxGrQNCn9bF0BUiXz5+HImOZXq1QOyWmyZh2pCrJ/yJkGlqTk
WYdDP+sBvyQS7N++bHbawq1mhrkwLoexlTtHJ6sCXmGntbWQHY5xN4M2wGZBed5FuIb8uzw/BxDj
dRD4qZwQT+xjVbyGiIEK8z5ihvFlI3zc+aQnr3XLW6x4qJo5wwn22zwzcv+jueFxIJyO3Gxpwb5N
uYAzYTqPMkk/FGF64k01GDW9RW43d2Fp1kxj4cxfD1/b6YUZmPAVjFOV6ReRfcuJkJxYSAMjKP4h
xzWr8M5l71JIJkUtO4VI3Eed4PIc57M+n9THImK2P7yF7WaW9r+PwfaN4mkS/CVQbAHr1aWqjVvU
CrCAuDO9dyVOBsj1zC5TOVe4TuPbB1L3IhI1QuBi/1Q22KP9j/XAO8xpmqK6ez/btY7Dxjjr57Et
zwMsCkFQZISr1ZXjGMnptLYcDUotI2329hpZwsXbbg+EpFo1BFeHVRzRzWkfZaotXxCbN3Wica+a
sDwa1i+RThs3HpuvsyEctdcsukjNaEdM3SxkmhZR9wcKCB1fYvEPKnZq1qWOdfSN4VM7JflVsqGZ
L8d6ExWB/rkGrGH8cDP3FUOdO4vBEj7NEdr0S73/6g7Uf3FnKfWaGgZ6XigKi487ulH9V2Z9soav
SKanfTA+fEFb/UYUR5INo5wl+O0X0BWPOvkJQ6y6TzNVX31itaDwsPqzgF1LpqFMrTYMAb//lDnR
ahAI5cxgIUS1fh9XN5sWBSPa8w+3b20HFpmwSg0cGH5LnLoLcbkEgrTKHas4qhGBq+N1lDTCef9y
Men7VSBjaRthmTlGnwFipz3VCYQPlQUz1T+hAX7oILM3K7B9KPC1DjW9QNJXUd7FFMKXNpmCLoDa
J8/WsJWCy+XBNajHg6LiITjb+ihjw3quLEBkBxpj2p36qCuanYjec2g+M/z/AZR3ZwZx70sAbu91
46kq4yZFFUgKCJWnHQHrsyfivpLP/F9tvkEdbsrhtRLrbjfA8dXh3gQhDVbzg0I+OGMwVX6lFDoN
Ooz6JB3G4iOY7OYL1tqMWHM2q9D/KSDVZ0xbDMh6cTiKjNaUfpGeBPVvGNZywGZ9iq9H8W20t/ov
JMJBhenAv3Y5Rf+ETQ1YNDorwhPeAjWCI255Gum/FBPcm2wpUgd4WGSPeXCfwlJsAUHRFoZGatRQ
4uO9CDRywiGMw2qv6PU6bx6gdpR5xyWEbcJr9tgff1NYmIoWIxnSP+44MambC9oOAFfNjGLqjH4k
0P3IRmmXwf/1nPoLZ3etMXA2MVqi0hWYCDNMj65CXIjWN7feODrSf5vrl0lHUQPIeMHuFv7GE/Z4
F/t+WmqVGRnsx9kecfjaRx9V+dWj1MD2EeLB1yki4nlBgGWi34oU9YY49obtKhp2fn87oiIa8fl2
AKoVGnOZk02aTo8UjqsoftTMLZtb1oqrDmARjxDTpb5j45gXdsS3TqlgVK7zT8EQkqP6T+f6Gkfz
di5MH/zvyMlJsOLdz+Mw4/cqLu0jODF871cRE10VzcmC07DD+0flTfWhJyZeZakocWpja0OaT6dC
lL5eWUhOcCcqtP/sbEv0eFznqGnJCAu8fm+isYJqtkwC7c8jVh0nu/Zdf7S37PqAV2ko/tF8+izQ
9OeQJbjNzCXKtMN1IyzAlRdJI3svH9e6aBLqBwQ0aO8MyeJOiOlOAp8YnmM3iGiaxd0MiwpK3O4e
p5LDU5QncxBKegBY6MybOeF9oUZLkDRlS2cB68lcuenPn0WRxFz5UOuE6H194o75AlvSah332R08
NthEP2DDjm6pWKUoxHzFy4Y4cbXn13cFxWbyw9DWhxI03pWTwg+x/SlX+v5SxcpNC5Zo5j4qkA8q
Riy3mrU55w0wlj9SPcmf7HZaR2+3SyhjRvlFe7yPSlBYjrByZPEce2p767fiPbqeSXpak3D4L8JN
UsYFV7n8QS/PjpqtVW4tnjwri6cCczawqPb0+rn2fNzYiuzPxtzmAhc6IkwRkg9iovdj7zLNX4GV
11a1WjjG60+FebmuwvSDD1a3YIQzPPS8D26XLlf4aa5BqSgMrMVkWyYOkVedqJTqZmL7a0faENyt
Yh1wRa7wTfbPMktShHg4KR7t/jx233ZTU0kXrxOjTCaGV8A0mvN5019mm42u8o33aYvxoDeLCajr
mpyUH37BMltEsscTcPxtq92N7DGoyVpb3jeXzx73mAOfTAzo3nGFDnQPvG70c2K45ZoUnNCVAnro
N5ex8TR5Tl1/031FTvqWTpbBQwOOvLh7uYmiAogNH2DGekVhunrUhrj1fibB+oWY7KNoHbt5BxZG
I5/hVwl4bMLcoQjLwAITH0RSEcgAXd1PAGOtJXRQXfcLVMVg2/cZmTMXcJv+ba/bgz04+Cz7KOjZ
uvNXwys6ipx511x/JBfH5cuG9sCVlq51rQ+A2LYmdEWtN16WDQ7KxYAvU+c4kW1ea86j9upM8IbO
7vz7K2t3+q1eoE8A/fqe7FhK3ali/bdlB58wMND+myNVkhyF/yaTwQ/7JPgzE0yEC4TMgkMP1Fzq
yOilW7v5dj+FGHh+wqXku0mtSRDlJS3Qr0BTjAvlYhhkNz+lu/5Vuy+ZPpFiOZOAzBwN2ORsFvGy
oi+ZreM9tlRxsDVWcZdBnqys2OO4CE7hwbTIqPOC6TAjoa5OEo1uveBLHbXcd/oedPJ0CQ4yypNl
Obt7Ol/BJg7NMkRcStLN99cFGNtuZYokZ+rE5Sc0NEUeOO4uc8/6MdTcmoTY0DDPo+lJHPJqX5IB
6A0Hx3FtnHliWAdj80ukN7iNrXaaPurFAPgg9/2DC64s4soaEu/e/pY3+xFR6+0tpvHB8EXmBB7u
RpZrqF3ZNx0OoINtQz6JwXu1oMRGUH2Qv4OMbIH3PZ4YeWWbzwMhhmCARbY3EVEDJrPVz3XwZIDi
GoMkLoVgyYF5jx97XW8+x7zfbg/Oezn5f9S1sv1saxyfddmoA9ZSvonCx3KJMyEzlVStiPPCvtQR
pF+W+GPyA83QVaLfXS96zW1MuKnjc78ukmDPsB/6h0Gw/b/cq6mJ7zu2e+YXe/kTnmgUGn36boXH
6MjXO/nm3I9UOLKPFa/8Bos5ae4ZGd+3fD3SydWOqIRqAUooRS+UwTC1OvIfcsawCCqeuf0wMIwn
VhscGdkKrKlo20YfAmGRxDWThgWffFY3Efr5JOQaTtbBZZU5/DR/0wIYugHNmm9CA2j6fENzT3lQ
JumfNyCTAiSDHO3vBEB8Ro/6Jj0CPd+YOSMfnSXh/A4n+NX6PnHcTYKo6T7fQV7Fv/ddiEL2rsC4
Y8Fjj/esNobED9nIwYojtYFI9K8NnnggbSfDlWT3JO2JbXg9pTg1bvQm0aaoIlhEXr7bx9UXSXiD
bgPtquxcfDPWnRYHq8h5gfBUw4e3oou21+HaFApy84S8oleze1WYEapCkvaoAKYYBFQR30gWT/bO
kYtBZAkM6lbr/I07RzRSpG+G4YsnUUXe9/6S9Gqk/l3p6B5C04ILTPoKDUxl/iOxQcHWXSikuTZQ
2Ye/1qLidCnFiq/ey6z+ab1mkMOyEjibN2j6yjjVzLl3t5Vm6dUxIHPUpha9q4YK//m7bbJykd6u
9g0ad2GqvTFRSSKATi3O0YZy556Zu0Vsh+++5YcMIUz51Xn6G3K8+laj3HoApwHPgaEaZlzwO3gE
eGxL8DrDmcMjrfOT/XnHab3xOLWRzKI+aF/Qf8YQCCELRHHaduQkYHej7k5Tw1lxh8uWRuTp9f9f
xkjBcKCNxiXwQpXi/2u+Rgy8xmEyI4jsAKMInDoBlFrTE0+29xw/jZbO038/WSHyJSk5QYt6eQjV
lmCuSYsGFgLdBMi7hSmlT1s3LMSf5DuBz5sDLqq5BIf9TKTsX02QQgA49k8D26GArRZ0TFKMxcqG
TKhQo8eH+S8q5v/F+jh2kmGxM1BBx8n4dGSmtr2yvn8GSlULFHD73ND9NNHdhfIzg8N4IPyt8c68
VcIeA2FhabHBUxq4Wirohc/C7UBZNGxC/stw+R7IzjXBqNDSyuR82DqEqjYa3W0fTG9N+Hzv7RQR
NDIE7ON4NlAHGDRru7KSHfxNTBo8M/gFfsRw02c2P8g+grFh3luI/wjGgmym0+0LN9juQscVkM07
Ln+yKpFpiyafb7aIUnUdSjHT4VDz6DbOleONKTyS2O1Jyqzt9idAlmKhclxDQPWaPf7SWgHNXRXV
Icy9YuCi0Zynttzu+SDb2sOPup4dDj+xe09Pd2cdxkiRG6rdB5VLynrnYkawAz4jnpLIBwGt7J3X
csXNjJlreXuZTy6tVFWTwm1CSZuZ58lpCnn/6j8VCVvcjPwQFyMAdUVfAzNVZW5qsputol+I3Ujy
CkkmLFEzo3VEfhHOYUyH5cpP5StRpY4yFmGhl928dmxDlAOFBIJ7b+eDn8FdyvmMvXY1jaLueO3f
eA1rYVah6HU9mSRMDXQvx/9o2J5zIPkm2S580SB7Zxul7l+WA4TYZv0J3HvGrqieVDwMMPWBznPc
IJx2f5J2EJmJncGaD0CM+dbYAfVsJbCVv8rgRuDD2lkTTsEJttTH0H4VRfqKS/OGV6gspNLabRLd
lz4zPD9rmcbXtQPwjZW+jnxRgW3/BVJa/GqGC/ZaZYt3VsZ2B0RTTu41fNnvp48St+EvIUiO3pu3
CUvEsqpeaFExVp89wRhxxN7cWJd5Ams0hi/U8fS5ryLwJq54yj/TLHf4vADtD1SqP/GCBX5BGpU1
M5rMIJSE5EmHeKxsgWzMtrWZhudOuPmW481kliASGv5puyan4+s2LJJSEq5EMUSkTNnHWvF5qXi/
nyr/GJV/Jl4D1ShkFIQuj1NVd6ev+Usc1cTmfhe1mF+KHTA7EEdvKe/x5baDRNK/Vo7VHPUPsTuO
bKr898wMHX6tphPx/HcgLVAWejt0ax3oaFs3xtt1Yn6jv5h941adt9WTe+8k8DfyzjeSxlbMveEd
qIFBAcZaXS1Kz0+8O8SDDGDMECZnYw/L+b123gGPwb7Kis5aMaJmsg3NIA6aNIySDNMkLJaQHRhL
ZK8ZlgIu52Yq7AaHQ4CpYhHke0cukgze1IIIpBtNDYIvHgVpaWtODCoXiOAQYwGoP6N2I8cX3TtU
YXmrGkTFSHxxDWJhUQCaZYSj2JIsH3oNPTqx2K2J7NTh4FDSO/vDR6hgiYH18QZSyRSAA/FBPciA
pHNA/CcqkjPMQ0huq+dcB6i/cfQIueTvihjf+0T9WI1ePnLuRUqdoCfCR+zEPY8+xt0nWn6Ojlrs
TgPfM6fHS5t9mX3W1y7U1wcdkIaGZpJ2NYyy8YbuO5BHIfgllAqahP6Gx0lpzV+I1eLL3RVG/L3G
fv/ORG402k5Zgew+ywnIyOGqACktm9F9Yrm3zcy5KeIIk58j1AqeFNdqDjn5OI7A/ZEkpccXiYQQ
Av06+A36REHr0TWCehl0TxJOdCXRD+3t6edZN0yTWhgEORRzfWxs2pL5FEJjJyY6kjBEZF4coF6M
ibYh2zZYzrbhahSAd6G1Sw7ML8z9Vm4hUD/hlcSr52/4LVeDj9GHqpaLK22A28byThRfmzkdPvGy
mCn1Q23GRgVk2XOonqPrDV3yXehAzrhIWznj+FjZwlIsnao8thlam5DAGQh3y1FlmXKkzq7q75jL
XS2SzJjb9fwEx45fw0EWeu7+cpG7e4fqukXKRs7aogapuPGqVBl77R3smYNGK+q6kGYdejspprGL
3aITzVJhsZthcfq1M0fxtsWS3wWRVIsVaqPvouE/4L78ix23UI19SVd7iComz+8Mfgxpsi9X2A6s
2SFVN4vRk9LHKa2EEb8YBtZakG3fg1TReJKQuuJVlmbGMGUcuM1qCYMXN7+8TZ80BOL/FCvu97j2
hUWZtShGVkzB8VHdl4s/7zSQtBmmHqo4vVIKMkXYmYh12jqAJwc1OW3x5pDyDOdlCSImdW3Y1MtA
97La2xer7tcxSs0lZNsh1uMChsTn64arQo1ykwKhTsjpHzar1bEfdNPgD0jzaBD0wXDQer5l3B8N
HNR9kTLwa+0DqngxWUcBQuieUITkwisgvNqriYAtUh4n2XxRUxKTbE1eF6bohsxqQEcKYAuXad/R
9x0Rnl/H19oaNAVURub/ZK9w5hpt3ah9Cs950iw+OSg/PqROU8tSudufslhiNUkKcPdLicS3pI5f
mSRsESLwdcWZ0LV5M6/2ZQxd087EAIm7qe0ZSNLREKDQp9O1B6DbcEXyw2H4Hf+gyKoHW9pyZcgE
ir3UzeznkaT6FBRW2vSP/clYwd4T9H+EM/eLRKTTD35QdfL/QjLw60PaY1gDg9APhxqttQlUl12W
8fR1QOiI9DnSODYc1tAkVKpyZfm7l0W1QtcHwW3GLGSh3ilxx23RbYM9SRtAZw5lCY4ZjeY42AvZ
o1ZTbxhfPOYVeJrGO85lk41svDH2vK0u9D3zrdrFR1YdEZvXKWgxbg6Lq8oCf3PR95JlnKrus4yt
tgj0ZJxh2Q30cmVjzmXDYg73ovBkPox9Rpqr8BE4aYXSPDeYOeU6vl564eLoox8OLms0iiM55xOr
3+XZlNAqRqgPwCwI52T6tOVLctc7vuHc08mrds8WTFFmSpfI+ZwzxVzeI+VB5E3EWJNWEW5VLYVV
VpIHaQ3rSqkwm5MJ1tbXcrzYUSKGRR8qLLUYiDomQwpA/rwNkVUlprFEdWvHEZlP6v6Z5XM8OG49
qAE+6ObiqmwNiSMAzRSrsT7wGiPAgN7NPoiVcFtjBGW0vjbo0+LsEOb9ZDANXyJkOGLRdvOgK2so
jSFYUscoslaeG5xVngkABTk+EDEXOor/3jnvVNfk6MrAe3z60au6VvOXP/dlRQI52pv7Rt5O9b05
W4jmk/8qN1HENBYL1aapmf4BKUqcCJkeFHJaPtU+MO7ZdYVcbtI/bLG8aNilnGFGCKCBwFt/N6zO
abe5XqiJSiUqAoHu98UW3HjMiXKEwy4lWCJQW4JJukLgiDcBx2MM5hibAoHQ/KjXHD6ldE4Flwbe
UmSKOGqpwTHCcR48Edq0701BmVKXrD4h8e5gCrDtUXG4M8dRSa+v5LPCbT7hVLAyk6B+eZM/qLUG
bB30Fc75VGYy15wWDLY4VlCnkWBuXUXjvFhjNo2z4sR/SSfZYz/8BAdJYLRUdFjxpDDO5CvrX0t7
8L/u7FjEZhIRsCcvpivQZNajsHO17jGm43qeZNd9nPZon5I3YCV0l+FTLTfoL3SfZ4vxo8qGfaA2
h286pK93O7BcwULyVf1RHBi74UL8Xd+ArdQ6t9VRrHAJWtB4PcGB2jAJ1ojgMsrgH9Cgobuf/kmj
ZUNjd/42zzpABwwC7w2yYPdYBE2JGrJ8pd2yfbsA0ZJ19h2POuFJhKglaGifsGiCptkywmHnhSqk
Clojw2Q8O4ktlIWB+2WY/ukpklQ/45QvYrdsi8RJXQ9SXFKm3b4b0qHIXvo5uthOtO3NtrebYQC+
Goc/Mh18a2xVFHXpDTUfjzS6qrv0RaVQpiji+g1DXmVX3d5tVwNYXHmwNuQLSZn4+YSsJ44ECTa8
WCVRtEoEIgiDR6iZLAF8d8yJfKdwOU0A6IGZphVT3F6DKcW4ED3BCWZUzzd02CwdFTfzd0fRS4i8
CCXjG0eIqRrJQMVimPh8f6DpeicfZ9vJnN7IAv7HXybpJI9UEckoKuSzvVe3WGr9wBL2CLRyF+xV
RWzQpa6ew/nuluCVDOId3Y8ztARn3ALycchLe+JzNSylssQMp/Py7QCJ8OI6gAcJuGxswEAdvMEf
4Vla5aoZuWiXRy0oIOnRtIeUWLawePsBwaBWpmgSugUKYklayyXnpjYIMx50mSpxhcXdBLY4FC5M
tWEKzIBSKfs7A8JDeHge1seD7UmH3LekeRXPs6/nfbG2YaJC/YQ4JWs489gLlNfv4Y7Yz5k7++g6
aHidnl8Hap3cJFqvRIBmdxghRxItfB0OBHC+1JOwmvj7ptNr3Oue7w6yhNHs41YFtjoWBON2haC9
Wfvl+d74YVz1leKxDyHT0kCH76+0Dime7adSEE74yO+EWU0Lca8/KneAg58Ff3MRce0lnaZ9LE+T
d7qL60tSePXuyOz+s7uKvgH4lOLjObZ8784OOW5RManEcQiMbo7+qM07XB9Pk+6zVAFEjqu362sU
4gT3B5TWKTzUocQQNxxGSDLFARSqafbNvgwxdqLmpoNhrR1lHc1uFHEWjmjR/JOT6kdUA2rFyw+s
kB3SVMeFppyMav/s5K0krJrSgKkKr2S1xdRXgOsFtu3V3TcMgOO6Uth/x0s1YI3c+gF6lkNGn3sF
8AAGrNAqwpz9s/9v+zqf5ZKx7JANy2rs03yEAPAtUBtdFURF1VeNu2c85oqR+iohNqnftJD08AfH
sL+pZq1cCcVHgqhiEeMyn0RCqSTwiiHiWlYLUjZ6n7rgDZQnI7Ka50cnPy7luZpYGkLUdorACmbN
uV4ldwMJtqh/i4e/BVDJ0nBO99aOq82QPObeww+CdIPQMqVsL+HP7+CCoWntKfcTYxixV3d41y5J
JH1totBUrVS/oEfwDce3NsRQXkDPp+5siqxhZ8D7rrBP3Rx0ZJihLVEgtNJoksSw/hmkMbTifBJI
rIGLg4THesaxAIBBJ55XHeDHetLjKerL5GlPz7qQOCsMnWB4lHnIgHBXd9U502UcTXaT2OIPt+Vi
NIkFsFrX7TPs4TbqY5PMlU+Oe4AOv7qjd0/Ohne+9UZZCoVWF5sqgZjt1eYzeS9EG6drbgJLeW0p
KlxxyQTN/QKkKz6qNcexNM3gaUcpJinq3LxDAZm3L/WC+wp77SuHYZzYU2FWLsNTrMV39JdlULq0
KGq+Jjjv6Q8pRdNqFerTu2+zGTgtgdGhIZXtdz+CPFuCb07okB4ViibC7ISMv73EfMpjTH8d9COO
T0rduZAKvBbVB8iEuT4D+8ns3f8R6aqTwBMl9ysPDUpak9P5imiUl7kKUxSNrQ/Z6afjt4f9Aidu
vTpVW4M/I+CBS99HukPF3Ri5wNFz94i0Ox/L21dz0k+FjH3nrlmXA2G4tgPsI9cDaWGuGTtuqe4B
wRkd1+GAB6rHRjkt1sdcOqzqMDbSTDB18paCQ81xwqDq8yH537InB8knqe5QCMlp020OxCApaL4A
iNDvuyyUIFi943qCz5tva/cYX+P2xo6/z/668RZ3TxHEmqbGqpU7ye5ncinwkeXBr8KFzrMOInBi
Z/EiG6df/QGSPwStKfUQntxWrPkujfr7hMSI0gGok5LSJ+o+8Y/Zp1CHMgT997sMYng6xNnVKj8L
5qnbekz85gr+h9eBC6AhWeF5T2hcPVqcddQZLqT08dweuM0tDMZDxcytPe3vy2pzl8wbZ9aRbLgB
OzFLmca3DXm8ZMa4ckR9pPzTwJSFXrvdOgZ9josk5wMnXr2z5oDx+NthSDenEEQpxl5hv9i3ZTE7
5rAap0TdAuyb3nmt4J7N420RfTAnVsz6D85IQFFgoUU8D3YQpZ0CKuAxR1vpo4oXrq+KwTn0J5A+
GgDRnEa+PZKfTnchOegZ4DHuPkqjMqO0lyvsqEo51/H5Dqof1xx+m80e2BhIl65oCNGjZ2ao5HCV
LWg/23pnZjuiKs/+fy2bNWVQdGHbsQRvvDSiEtn9dkSw83GwniAg6qbtpQ2DhB0NdHUVUqEtvViO
j7J+3tYaLPXaoEz+ubr5vsdFBubR6uNS+0U5L+8Dhqft/zAvJipJFNGebP22Bpi/jYx5x+H2/Ci6
Bvb3O//0DKnn0GIzLCrsPIsEklEIGevfJgBRJhXTBo2wEPgQhlycXIZlMA4pmd6NhOmhDXdN72lA
Y5z0mNU7NbZ1ovq6ab6wADSziniu8ifHB8CLIZJH3OJAAb/K9EehQ+gOZ1wMq5z6VPNWgO64LYG8
Iwwc8xCAFNymWQsYdaBiB1/4ngiSyCMBfI5yU128oWy/NlAsTOjVdmMSpkXYwOG9VWfxeH8/1VQ3
HDXdF6lijhAkCLu+v/TIrdzGiyLLlaB2gFPghLVB5HiJOCsaedYv+91xDKYeXA/efIUwTg3nW2CU
qXgb72cRptfmJN4XEOxCP52EshFi1E51WBxL/xBG6iDkdI7uli00ISxP9hgpFpEc2M5LQAIYwT3k
A4ZTH+RLTh5cVCXtiL2vChUkWp5vHKW/ZCNJzHAo1RqezijEeo3cwF+2ImrV6dXv2r+zhu/uXo8s
rqgfR2orweffQZFKxdue4j1Xl4Ahr+IC+zZLYfJKMh203xd2Qg2xFh5T735IO+WcCQIJBaoGxC99
DpZObWcNIX5L3gGy8oYzyIBwRSGvDONfN0g5IAyFMxN6OSvyzF3csiL7mriz3j3tB0F/MyLhMPf+
z+sHf2o91NZ2fv5jv4gIX7SrOMvIiUo7wU54RsQ09vwMFO5FoA6wtch2mTm58zZmUefH5VirxoMK
enlaevFv5xMJ+hq0AuEO2LJqsFrw+DuvpJDQr3s+9VNR3WyUxa1NLsQtc6+oyzYJbPN27eOariPB
s8Zq8NOv6zRQqjVdm5gZluvlk2TQSxsjQEAK/Rq6qNs+DVA2Ceel2HqvBktkUyseRRuGm7xgZoR3
PP4aL9gWFDeQaqnkG7lQ8/LOovCR5Eb65mrK+r3vNsdb1EGFlHycRk7Vw6ccj71LsjYKI2Et3h2D
zCQEKH1ELJkd07Mf5SOInuGtPaZZOIRuJVQHztKzuGQWqD5x2kKcUBGh2ml9a2mG/NeLbNqTAldC
d4G2VdPpGGGoADc+m9bcrMxjB3LLtTev1gdAq1bSY08G/sh3G+Ar1hm18lIzuZR1J/zym2Z7kfIW
q+HuD6/TWxyCaoDu1RlDuihd0Mp/PbshuNPl2mJqROUBKtLmfv6HSOl2Z1KiBUCSc1OwU8FoNb1Z
jNHoS313C/X8EeSlSSdYtrrwk+5se0zuM9mzqDZnbOMHcaF4EosFCvybJQDpJNXW3yFXN9CnkpIt
voLw/s0gFlcy0L9TCvsSwHkTS/D340H2sX8nW3OIVhf4Unozr/FpFP6l0bJsCVHcTyPz4q6P8+xx
K5gvalZupkjXBKvMUluMqFFp0yLQu7tsHwWGumLs8p78q2LrqzOeUuEd0Uxl+ueuHh3QQ56TW4/v
836g1nmah8AeVRJ1piyQVebRUs5i2YW2MnZX5NzeyPSLWkYiv3ATQK0fm1caXX5NIRiv8v/dC0Td
LUKN3wgH5aHm4cM/vrA9sAofOKYhzNL2xMai+8R/JQmHtaJgWPc54qi0cqA3DLudZEEdJ+DP2aJ0
xC6XA3AXeg0jgSsuMmblCwY1aDvT8VQmXHjJhsrOZfsqbyXuYDOcCfEROxoGuIunhRJc7xc7zHzy
j/p2/ITiwW5kW1vJfvdFInUH34VFqmbS0K/Q3WHkYP5i/eeItOFWlOaTClhuO+ho6lyGqtv2bQ9W
Bh/Z3ocKyiYyWb2C1kVJcA2Anniq70LBr68szgjx/Jb+t60ZqA2lSQcsXiuu14c99kxtxBn74en6
8p8pROkzfKodrXGqA5HlEcbB/ikt5QuHCXVcvSsxJmkeG06+Es+ysalq1PiFpLlEtzUrtR8HG8RP
0vm89YpYjfna5N6ISGYjRcNr+9F+9Gt5J8y13P0gkBoaRZvFUwwpm28vHRVxv32a5QFBsO/GpkXc
uR/qOlCiqeQuvtQI5N7WWyZlHpMiTMdlf0GdwJH3hYvBLu7YuGW8YsWuqq/WuYPmWF4wlI0L5R7k
v8m6q81UwkuvENUvPbwyIcLUcJQed5wVR6ugscqoqMYPGpkx/zPAZX3Ni+ZzU7gYacKZDosSDYeR
AnYNVmCA57kvXC7z68qjWtHFPQmrWBLjJXmx994lBCykb6seqcG66QRBCojwTpP0+Dz6hhwOHanh
dNPSdIU/KQYuMKo0TysKu+qloaf0CLkXGsy6ZGQydNfNL4oLvCX8bbb7L8KqiHzKgLpYiYpSP5LV
gkdR7cYVn1HoD+Fb1BBtMKHt1LK6eDEIqjdMBHg1UlYKqYarEnm/VpXIHvS5OKDIYupAXu8wlqeu
9XSLsWVhaDXOeWh3Bxyss3uU+quJNUjNI0zD2PoXzjMUThV8PKN+27/tpNGlfA2I+dhsbIbvXnn/
A/Kb2S4Koc59A8CkWru9znayj6mC0RKZEcif9VXirO7f6V/h0mt6mSlaNnb8teNNTGjaav/4Zjiz
NscuUM5USvjbIJtuDrE0I6qwYT1NKmXS7qgeituDbsy+xNx7Gb+F0zwC7vylE0c6RiOg7jZzq55x
v7JqvqERNOthsC3FvjNGrdmhioCxq9ZbEXLYWZ8l5nsY5TAWOWGLofYuYKCxqL5HT76ErHkWsiiO
8rjHockRgnVVTgrhBSzIEV/Sf9ZjH8+06+e0gsvPVPb+NbraqvahSYBdqILjPapp1u2MaiCi7Lah
4QA7qajBAft63H2SF6x3K41ufxbbvN9P5+tY36ZJ8eRSICsNXnh14NdpRq2BbaDlorzhfrKypmi9
a2TgBczlWyMdiwFcBbt54LyUFU17e47jia0UJohfxi7Ha1hbCB8jLRGNNg4a6aiI14yFCnhVWUFC
l7hUJkJENTK8CPgscU5omGUISCoGFWSErgqSPdpjFlI63kXe1HF1QDCXZmbx8n17x+CxK7aruUXq
U9cWttTl3LyPDvpoIqGwHKq5PCSFURPfmeXPxUkVn/f4lb7swdVRECivmIMbrhs1OHlkr3P7xA1G
95Ya9NY/faPba32N/MP7sde6iWCx28enhCGYRCnIMiSLtmsLvwXqVJiYJLJIVTYLs3X1paSq3sGk
tnffobFd/mBqyBpfYQq8VZr/R9JnvkOf0hX9p8NccIYlqAeiL3nP+mHbC9U71zK8H5I4cEWZPtZA
VfxsNd7DKClA4sz6P8agTw27Aafx2xsTS7cqPkGQpZy8D74VJvbxu7wRRisWvI00OPNxSJPWr7yM
g39ZBNR97wPP8rvelUugTFm65VU00EGeymw3LfcRqPBWXd2ILTqweHdj90Rx7FqjSrFDnnCvwGmy
7qLUi8MsizVHoRu1HfGDyYgrHic5deU8rv1nQoR0Rod6WC/jwiiHUsafqApyFMtxBo6dONgs+3zT
tI4hgsdfgGP9rIB1zo1jzdpUTBwXaDFvFcpT1MZgGLTKZWwxPO/AW/3ez/B1tF9ev0NC26JEfPMz
/oUnAnnnk07a7NE+ObxeP53D7COR5AOdIQR0x0LRXOGshi5zyJ3wWZpPUJjgYEzV1XU344dtpbv3
9U0GB5V3I9X4Pz2+oT9pWhxLbWHOLqYlBJZq18vBTsUuqSQ7mclAvOmMj5Hv2kvHajnPHCfUR8/n
xnAEc4Ui3DizDYQgUvBwokS3LtpVCQ5fZjSWisrPbdQYjES7PjBK9jiSy4A7TRFurEOAqbe/oTxO
DXd6ZQ/MVlTOht1Xp+QQ/TgzU8V1lpOv9qy86g/2UamfRkfNTx8uZqTEzt6sq3eyxYOCQFu09kbZ
Ilefdzs2iUfm2psa9KCcU5nv89fYSn0SbCVQ8eHOldPaH4XA5EdZjOW3Qj2/KuKStfG6dwkBRx2M
ymoewVbijZpAoPG3emlMHZz13qoOYmU3qNE2lTEIPNKAxFc+c0+G4paP58st8FUhJZBOkWdOnRxi
Zh/dh5QLBOT3bYJD2I5QeYoyXx4E0q3IThsnu62E1oB8XE7/qfSN2Lv4DeAzKSGNBIvloV9/MYYv
i+plL++iCLdF9fktbS7nKIq4vsYRgPEY/UUlfMdZdjkCubZGqKYLC/hTk4QG8oeWQnPMixx0SsNQ
oDpGO9bVxJSteY0hkCt+ZjThffNW7tQKN8hx8AOgeSxLnMz1lXv8+f4QXGulBI8X0yqNQvVxf9nd
6xoYw64qZQRcLS6IC2U5+7etxOxAhuDkvD7HQrMQEzvRxH6J6ME6J4nWCfUrM3Eh7UUcIuFVKjQG
wP9dWujnj1/lOY9tPI+ev3jdNVI/4ffWhqwYfrWU3LhIQfWyXwMCdk46DLhi1cZm5TKx78freGtH
TZDp/wyOT9PsgCT0YPAkOkck9PF3ioB0L6rpCTbvObRqPWfTt0Uc7zcKyKlb3WqqjFWE1IzyePhx
kqvvJO6t5/ANHjz0QmF36/jGHN8D9zB01+AooKek0jovPlApj3GyIXh5quz6Gw1GsFUz9Hq01fdE
r6Lo5UtYYiKMILOrnNss3W4NcJVOzMrB1b/9IuzbSJPi59pDViax97gHcutOPZnQ4+fMP5sn63AI
eFB6ZdBcgP1tsBqCRsizMLUcI/Waa2UuyBt0WOC3JXg/W63mTGNme5V9XpCEzLSCLeppzCHnXzqO
F4Y5YzWrI5eCbTJMmMIAc4m5cQrFu+dnEzL9xR/5ZYAbSYJmcuYgXCnP+rACYMmaUw9LLcMyNyfU
3lbLY9xLmfUZPtc0AHaYWDMZ0vlz80JGkLjZnw080V8k0JujAaN1cZ9I/jJVZ0JySahQd4yprTZo
/vKaHF5VoSTwWi6CPUKToxg0FUgoVQ2soZiGCQF1GMWb8Nayvoa4BNcmrY58hFyxMx/T5v32n604
YT7t2p8vCfaQTMARGgZEXLraGHOJN7qzZ1rOCgGzWJ0py4qnt+v7qAhEp1+5ZghTZIqNzqpT5ahL
mbZbgz3Xp+qvPxjbmXl6VSwXgxevtaiiZYQ6ELDxWUshbcwlqUhsZQKhdgVIuuJyaxrGwl3ExHXV
Hz9cw4dmHILrbcjmWrlrTLXGTKJbGhkT3I5qF1CfaG++i4uWmNp3CacBS5GIbziMULl4PnilnM1z
0EoKgJUklFIJS0ETQOfwtlguOeubjliHg2ffXpf0x6h1llnwyvowWSWWR8HcH4kvbBlZihFyKYEY
wSAhPAGamdIl+MGkj8jEz7oPaN7nlbXqRblGTLuuwslPYfQu19F8V8hmNpVfgj2cLv6jvVgWMTOb
R/MZXc1aKdU8nVWmuJy77IcsvTm5NcY590l+gpYI1J6T4FFu/tL0Iyt6Pl0FIU7PfVm4M64v67PI
DtCPOSCDM3aFZutd1IIJ+WyUo8tt81GahllcsHuKbqHtW+mDyR+6q7FtLg3g2ivxHTjbR2IYWx1l
b2Lh0UehcCoxUeZ+uugtr9JolR5t6sMi2RYEeogmDu7JmLv3xYow79ti28Sl81vEuadTi50thnju
ttvASNZOFiDgLGe6mmeDq4IGUJ1NxS56uXQ1tvwsnTVwoT2Sy9buP25dLy0XAN6TLTxyGrdeyvMo
iYumy0gx/WvhgonoxGWKxk1tTuahfA2M7oXBMdRgu77H/298s1XAA7TeovtOmRQRdRRVcWQzf4/3
PUoRPwrM0wh2RcoDMCx70kDGNWrNQcdegeL4RWlqN7S5E41bCUmP+/RaxV96S/GTSqjibiew0LGA
rRSv4FVzljd2OD77IPJVqCQpfHB1D3HCxgD7V2HuQFpmQDxiwB1nAKFZ4DzP0fsBV1Sjrfu9rMqv
SsFH5rJc/65GkW4vshhXicOmaK+msYDdv8J6m/BZl9m9afQTuzcDNS1psO6GSLD2DbD/qoDOvAmH
mob6ToB6uBP0XIhnTSb9C6xeJUZJW9XP+dLq39Qi3kyqrBWGLF53F0vBHLLRqN0IAgk+gs5Dpe5I
IweiEJ4/Ww/oWoFfiVt6YmjuzggYZqx9zGozneWW5bEe74rR484qmQc+H7k6xMP9lepxdr81lAIL
a+zs8XCjwuJodFvkgwHt+WPB5Y78bKtyuPg2H8cD86p8H0+DSfsZCElHjoP/RTovJe11SId/cBHZ
UOQRNijI2l25+sFKCKU5uqCFTs4BLe719ejll2pXWgd0I59PSKDMnA2YEI/sMrAUWpvpuTtdQlPF
6/e4UQKzvXoxogW78whwqpMDeAas9I5L70C1sA6Ntm6iWYcIixMctfvKA+CvqwN7iIlwhWHR6ibt
gkBzVjV/BW4duP0tiZSgT3rRaJu9SdTsW9WIrksmlDeKqLSJUhTtBKRkDqRvccEhYQ4IEBLxJyNK
64C6HLaofpA08T2JJRM5SHrrwqRHw987WcZSVGZFtk17UoGP7SBMPYCp3QmyRiVLn+X1SnqkEtmW
3XO3R+zHGJQIrLtiZmXuP15uulBPu/WdFHMZe28cKIRP86jHCRK0o+CGh4LCSD2kHivn8gyjMlH4
+/lyivu2LRUi/bJqICyrtcigiCULPGhp53LPHrKlZgSa2Vu1pFUHZIBRuAazxNdiCHr3d2tbswHp
5yuCBTTyeHs2suZBfupeO2vvwYZkMb6PqA0F94Cvb8YKwa/TXp5ix+Vua6igyINz5Mi/GNm06lsv
R0AFjphb56EpIz8q+1sPJCOoDP/zob7QRiRmRNsln1Gnec9erPSxC/cAZpY4DMc3FfvFMbNI8Cjo
RiwsdHud42xQzzg/FZTKe9z7EoWjCRQOBmflcK1HqVUP2a48ip5XpKNu/U+sMvGnF+LlC03ycbj3
hAFt+Bc6STZRBIwNctH8IkK0e5a6uY3BIQzDsZUON6mBx+5NnPFuX3McZKBuKgpkR5ZOHTHVUtCH
RuQ9Lhf02GERRRrtZX8qnXAye+56WS4zZ79qSWQj4ZBOc+oxiEo4tHCyr0BgiKxbM9GmU3SAHlqN
bp2Y9aT9d4NXGCkt+QKRggXV9qClmmvMAY77pLsRR7ajdqZYQGWURTeugB5xeqKhr4uoNhviXtT0
SSer8cdcKtWxMHRDCqUsjIozgHrwmqivOslBpX1CfaDRIAGTHmrjMmrQ2BqFPeIXTkF+eiyC8jhJ
k4lcTyN/y82bdUvWGpdma+ChnTZJztFWHTa0aJJKbdNY+mxnaP5KYKpEUej3OA3sGoCfRGoiVze/
SsMl6GuO9A0PSriciX1x6fXNdvoUTVbsYPtOaHIdzITl2Tj8V03UnQ/8vGZ0aTdcTpJ7as+lxQ0A
juD9SQqmWtQIyKsa4HWFrdQ0VIqOXY8rBluuZCGFnnCAosqL2Dte9IaUYd6FimP+2+mQo20i0mrc
Cl8rYzbfq/YgNT0hIaDk/J6KtbIr0QqhtVLTgcgZi6c7XVkY4eAcSWAxz01YiXGo9eSYBYwdOBSF
jxgX9fdPPsyFBlO3/eQriWctxGoA4wzR/5TLuKZqhnBATcN5Q84/7UbEM00uVzHunU0gmJN/RqcT
L44U6fG6IhUoGOFw5HnplTDZXhFHUmG/z5ExZe4/3Y2T5Q2QbWVzHw+S7jd51vUmXi9XHBPSX7ig
m2Hzj7GJLiyasIB8jFbAL7rDGxJjSdDsyFvBOHOG2wENZp4ySZiE8Q1uqevS1o1EJqtshTMW76Xp
0tQ0MCd7Qo6yxORsQ6E0PWr7M638kINKYECZzxNHPpAmF9m3CsWve/76+W7KNXGpLFdhdLZkGtlV
6+4kMhVrV8aCrCJjHrTM064xXkqiUsvkxHdQcs35g+ThLAwUQlunvo1NQNtbmzjADUMzAOtGIWso
AtVa+a1ForHaYyFu+kS7KUJLZJw9W1l8lJhb4W0aJrutUtl2vqQMN+SyKI49ePNaMgR65EquJ++8
pbE05JxtJydzZxJRYfy3p7n+53TI4TTXs1m6K1Sxpfg3ZomAaqik6fH0+6OjF7WSQkgi4ow5mlQe
iegalyHS902MgmkE/mUvU1X5AooZVHyQknMYf0mPjBbaK2yIowrYY7mcWraeKH6mCotvqbfZoLSF
Z0wYREkat7AhDIUdH3ZxbSOffAHcOtyw5YoVsw3TjitBAl+4ZOfMD94+MiMX+sc6ZNOA9hzbkAle
vXZr6bqW/WaVYJuGINHL58ZZ3ZWBawtimx4//jpDHA60/DswHLbAU2KCelVVKy4wty2QitYXxF/R
DxauooYlc0W2fU5xKebvAeObut9sNnGwKiQvgGjSGbQWMZBJg44fDQm9qGxMcWsNtr8rmTg9aMiY
zKPLRjJNwvhBuIC+R0vL+SQr6O/JpzwqVdpo+2C7KDdgdHgLBxjADztTYNmpssmx58SXrJhUi8VJ
R6f/Ri8f8wMsnXM2MMIK7ChzrCs/7cgY91XlGqfB7tzz5XaXte4muaZYs0eMggAZn5hmQyU+mdEK
MgvuXINfG0Vz/3+vUX5rnaDOCquXOgYg2tuFNxniq87FnUHw7slKvkLlf26nKxifeVD/LKJJnZsQ
+v7ki5sqZUJfY1EWYDyhkW8JyCag2FxyprCB6goZSNyarKHTWtqzYEQe8owj5y2HsIp/X7HGM4gg
ChImh1/NnSSWakVeqyagdFxN0Ti0hT3WRQGDGbfu48m+6+TZWGGDuwatZ8E28YeSBjs8eesJdMRT
00VBGTn8MxXvmh2OrL3grJhTtPxyR84uGwRqOQPcrmiLN8y4pWM/SE8D8yrEwN2hXjZ0FAajFtUj
lRCXR+PUzzd1CNDih6JUmjnmkNzQ/jAQ8zE71U50pXlzMpCu0h4/RZl6hzvazf0RQTGfhQjsj7i9
KN87uj7VMBBFsefYllss1fHvdzo+sH0yN3WLBHF52+pU5gLHeimfDPGvWFRbgSkZPmACQ9JivcUP
X8A6qnEp3lIH0HwU4EDHe53fiD3UY1q9UBvJXIopBHhgmsPy0LMedkOMDz589rsvvgXGmqWQx6Fq
7r8CzWagzo1ENgFj9sSGvpUkjE2qVoytmaL/SWIqAaCpxPij3itXGZV+WFCNVKSE7qkThURuYJu1
OuVg1UyuT16A3+f8QS7EcW5782tZ/+0O4T1ib5Bx/oKMkCR3Us2dxdGnBEyXXG9Pfo7BBhDBDkX3
E+3OSnzqQSyoG519sglouvffNzZ6NsUA8AcPm5WxVA1yXCAgg//XYMcf6Hxd+Nygd/0OCgZi3ekl
7wyCdChRyVc6qIkF9j7Hjart6AtYHjg3Elez467nVYk6GMxjD4DP/BsfM3Y6BLHOgR6EubpMmOWt
0/OJfYDJgfOKSs8FbfM+v0G913SIg87izV4d8Wyytn3hYwn598+xpQz600ZMhURKFC915DAKlhYV
4X+WZJ2rQ56yPazkmMGMUtptguclWjBT+5K/EZgtWf396zWmOfd2pRMKSH1EegddqAcyUQ6KwBlE
wBuhBnpx0y6tAcQMfnDbY0SzQK5yVR7a8Y7muymSVvx4uDg34o4XRlWCVgVTvuUJLQM7pU0S+t3K
v9oZCf1AEmbZjgJ+LlscBcOVNg39EM/OndZlqzdstvxLybTvGWGqkC+ZchMQzr1TOi1SczPIMJsR
1JS2N9hfmfyIjcy2P/n7Vm1xA4zI5lmflubfhepjJbQKBcyz8V+wIevikxxh5MZX6bEFS15pCAHD
nRg5ziMXa2uSmsC9cg/GIQK5JU5UxWkDFo7dYyycMQ0YZ9ifwNhs8thwjshFdR2ySjatz4TNvnL7
OmqObPjBKE4y6y5bcNCAL4+p8BVAIjzp4ltZJT8oyzBX6h0NNQi5NGGubie3ZOeY9WtXMvmQMZ42
Lg8IPpv6/HtxiGlb1vSKFI1XcmCAbbhccJTav6NOfKBBQ7LvXW0msaAs8dIziU/fO9tIPxU8i6Go
++qRrf1wIew3jG3e3OHqMUZYG9GCDbg21Af1sb4R+xQXnewUopggJkkXBaVWljfncmvHru4dsSxn
86HbikTPduhLlfhICSjKM6lAeRlRaDRJRbI1BqSBeJUEER8fml/qN6YA6Wxl5RDXbu8IUe4ewwRr